module BrCondArea( // @[:@3.2]
  input  [31:0] io_rs1, // @[:@6.4]
  input  [31:0] io_rs2, // @[:@6.4]
  input  [2:0]  io_br_type, // @[:@6.4]
  output        io_taken // @[:@6.4]
);
  wire [32:0] _T_13; // @[BrCond.scala 37:21:@8.4]
  wire [32:0] _T_14; // @[BrCond.scala 37:21:@9.4]
  wire [31:0] diff; // @[BrCond.scala 37:21:@10.4]
  wire  neq; // @[BrCond.scala 38:19:@11.4]
  wire  eq; // @[BrCond.scala 39:14:@12.4]
  wire  _T_17; // @[BrCond.scala 40:26:@13.4]
  wire  _T_18; // @[BrCond.scala 40:45:@14.4]
  wire  isSameSign; // @[BrCond.scala 40:35:@15.4]
  wire  _T_19; // @[BrCond.scala 41:34:@16.4]
  wire  lt; // @[BrCond.scala 41:17:@18.4]
  wire  ltu; // @[BrCond.scala 42:17:@21.4]
  wire  ge; // @[BrCond.scala 43:14:@22.4]
  wire  geu; // @[BrCond.scala 44:14:@23.4]
  wire  _T_78; // @[BrCond.scala 46:18:@24.4]
  wire  _T_79; // @[BrCond.scala 46:29:@25.4]
  wire  _T_80; // @[BrCond.scala 47:18:@26.4]
  wire  _T_81; // @[BrCond.scala 47:29:@27.4]
  wire  _T_82; // @[BrCond.scala 46:36:@28.4]
  wire  _T_83; // @[BrCond.scala 48:18:@29.4]
  wire  _T_84; // @[BrCond.scala 48:29:@30.4]
  wire  _T_85; // @[BrCond.scala 47:37:@31.4]
  wire  _T_86; // @[BrCond.scala 49:18:@32.4]
  wire  _T_87; // @[BrCond.scala 49:29:@33.4]
  wire  _T_88; // @[BrCond.scala 48:36:@34.4]
  wire  _T_89; // @[BrCond.scala 50:18:@35.4]
  wire  _T_90; // @[BrCond.scala 50:30:@36.4]
  wire  _T_91; // @[BrCond.scala 49:36:@37.4]
  wire  _T_92; // @[BrCond.scala 51:18:@38.4]
  wire  _T_93; // @[BrCond.scala 51:30:@39.4]
  wire  _T_94; // @[BrCond.scala 50:38:@40.4]
  assign _T_13 = io_rs1 - io_rs2; // @[BrCond.scala 37:21:@8.4]
  assign _T_14 = $unsigned(_T_13); // @[BrCond.scala 37:21:@9.4]
  assign diff = _T_14[31:0]; // @[BrCond.scala 37:21:@10.4]
  assign neq = diff != 32'h0; // @[BrCond.scala 38:19:@11.4]
  assign eq = neq == 1'h0; // @[BrCond.scala 39:14:@12.4]
  assign _T_17 = io_rs1[31]; // @[BrCond.scala 40:26:@13.4]
  assign _T_18 = io_rs2[31]; // @[BrCond.scala 40:45:@14.4]
  assign isSameSign = _T_17 == _T_18; // @[BrCond.scala 40:35:@15.4]
  assign _T_19 = diff[31]; // @[BrCond.scala 41:34:@16.4]
  assign lt = isSameSign ? _T_19 : _T_17; // @[BrCond.scala 41:17:@18.4]
  assign ltu = isSameSign ? _T_19 : _T_18; // @[BrCond.scala 42:17:@21.4]
  assign ge = lt == 1'h0; // @[BrCond.scala 43:14:@22.4]
  assign geu = ltu == 1'h0; // @[BrCond.scala 44:14:@23.4]
  assign _T_78 = io_br_type == 3'h3; // @[BrCond.scala 46:18:@24.4]
  assign _T_79 = _T_78 & eq; // @[BrCond.scala 46:29:@25.4]
  assign _T_80 = io_br_type == 3'h6; // @[BrCond.scala 47:18:@26.4]
  assign _T_81 = _T_80 & neq; // @[BrCond.scala 47:29:@27.4]
  assign _T_82 = _T_79 | _T_81; // @[BrCond.scala 46:36:@28.4]
  assign _T_83 = io_br_type == 3'h2; // @[BrCond.scala 48:18:@29.4]
  assign _T_84 = _T_83 & lt; // @[BrCond.scala 48:29:@30.4]
  assign _T_85 = _T_82 | _T_84; // @[BrCond.scala 47:37:@31.4]
  assign _T_86 = io_br_type == 3'h5; // @[BrCond.scala 49:18:@32.4]
  assign _T_87 = _T_86 & ge; // @[BrCond.scala 49:29:@33.4]
  assign _T_88 = _T_85 | _T_87; // @[BrCond.scala 48:36:@34.4]
  assign _T_89 = io_br_type == 3'h1; // @[BrCond.scala 50:18:@35.4]
  assign _T_90 = _T_89 & ltu; // @[BrCond.scala 50:30:@36.4]
  assign _T_91 = _T_88 | _T_90; // @[BrCond.scala 49:36:@37.4]
  assign _T_92 = io_br_type == 3'h4; // @[BrCond.scala 51:18:@38.4]
  assign _T_93 = _T_92 & geu; // @[BrCond.scala 51:30:@39.4]
  assign _T_94 = _T_91 | _T_93; // @[BrCond.scala 50:38:@40.4]
  assign io_taken = _T_94;
endmodule
module Control( // @[:@43.2]
  input  [31:0] io_inst, // @[:@46.4]
  output [2:0]  io_br_type // @[:@46.4]
);
  wire [31:0] _T_35; // @[Lookup.scala 9:38:@48.4]
  wire  _T_36; // @[Lookup.scala 9:38:@49.4]
  wire  _T_40; // @[Lookup.scala 9:38:@51.4]
  wire  _T_44; // @[Lookup.scala 9:38:@53.4]
  wire [31:0] _T_47; // @[Lookup.scala 9:38:@54.4]
  wire  _T_48; // @[Lookup.scala 9:38:@55.4]
  wire  _T_52; // @[Lookup.scala 9:38:@57.4]
  wire  _T_56; // @[Lookup.scala 9:38:@59.4]
  wire  _T_60; // @[Lookup.scala 9:38:@61.4]
  wire  _T_64; // @[Lookup.scala 9:38:@63.4]
  wire  _T_68; // @[Lookup.scala 9:38:@65.4]
  wire  _T_72; // @[Lookup.scala 9:38:@67.4]
  wire [2:0] _T_508; // @[Lookup.scala 11:37:@430.4]
  wire [2:0] _T_509; // @[Lookup.scala 11:37:@431.4]
  wire [2:0] _T_510; // @[Lookup.scala 11:37:@432.4]
  wire [2:0] _T_511; // @[Lookup.scala 11:37:@433.4]
  wire [2:0] _T_512; // @[Lookup.scala 11:37:@434.4]
  wire [2:0] _T_513; // @[Lookup.scala 11:37:@435.4]
  wire [2:0] _T_514; // @[Lookup.scala 11:37:@436.4]
  wire [2:0] _T_515; // @[Lookup.scala 11:37:@437.4]
  wire [2:0] _T_516; // @[Lookup.scala 11:37:@438.4]
  wire [2:0] ctrlSignals_5; // @[Lookup.scala 11:37:@439.4]
  assign _T_35 = io_inst & 32'h7f; // @[Lookup.scala 9:38:@48.4]
  assign _T_36 = 32'h37 == _T_35; // @[Lookup.scala 9:38:@49.4]
  assign _T_40 = 32'h17 == _T_35; // @[Lookup.scala 9:38:@51.4]
  assign _T_44 = 32'h6f == _T_35; // @[Lookup.scala 9:38:@53.4]
  assign _T_47 = io_inst & 32'h707f; // @[Lookup.scala 9:38:@54.4]
  assign _T_48 = 32'h67 == _T_47; // @[Lookup.scala 9:38:@55.4]
  assign _T_52 = 32'h63 == _T_47; // @[Lookup.scala 9:38:@57.4]
  assign _T_56 = 32'h1063 == _T_47; // @[Lookup.scala 9:38:@59.4]
  assign _T_60 = 32'h4063 == _T_47; // @[Lookup.scala 9:38:@61.4]
  assign _T_64 = 32'h5063 == _T_47; // @[Lookup.scala 9:38:@63.4]
  assign _T_68 = 32'h6063 == _T_47; // @[Lookup.scala 9:38:@65.4]
  assign _T_72 = 32'h7063 == _T_47; // @[Lookup.scala 9:38:@67.4]
  assign _T_508 = _T_72 ? 3'h4 : 3'h0; // @[Lookup.scala 11:37:@430.4]
  assign _T_509 = _T_68 ? 3'h1 : _T_508; // @[Lookup.scala 11:37:@431.4]
  assign _T_510 = _T_64 ? 3'h5 : _T_509; // @[Lookup.scala 11:37:@432.4]
  assign _T_511 = _T_60 ? 3'h2 : _T_510; // @[Lookup.scala 11:37:@433.4]
  assign _T_512 = _T_56 ? 3'h6 : _T_511; // @[Lookup.scala 11:37:@434.4]
  assign _T_513 = _T_52 ? 3'h3 : _T_512; // @[Lookup.scala 11:37:@435.4]
  assign _T_514 = _T_48 ? 3'h0 : _T_513; // @[Lookup.scala 11:37:@436.4]
  assign _T_515 = _T_44 ? 3'h0 : _T_514; // @[Lookup.scala 11:37:@437.4]
  assign _T_516 = _T_40 ? 3'h0 : _T_515; // @[Lookup.scala 11:37:@438.4]
  assign ctrlSignals_5 = _T_36 ? 3'h0 : _T_516; // @[Lookup.scala 11:37:@439.4]
  assign io_br_type = ctrlSignals_5;
endmodule
module BrCondTester( // @[:@799.2]
  input   clock, // @[:@800.4]
  input   reset // @[:@801.4]
);
  wire [31:0] dut_io_rs1; // @[BrCondTests.scala 11:19:@804.4]
  wire [31:0] dut_io_rs2; // @[BrCondTests.scala 11:19:@804.4]
  wire [2:0] dut_io_br_type; // @[BrCondTests.scala 11:19:@804.4]
  wire  dut_io_taken; // @[BrCondTests.scala 11:19:@804.4]
  wire [31:0] ctrl_io_inst; // @[BrCondTests.scala 12:20:@807.4]
  wire [2:0] ctrl_io_br_type; // @[BrCondTests.scala 12:20:@807.4]
  reg [5:0] value; // @[Counter.scala 26:33:@810.4]
  reg [31:0] _RAND_0;
  wire  done; // @[Counter.scala 34:24:@812.6]
  wire [6:0] _T_1618; // @[Counter.scala 35:22:@813.6]
  wire [5:0] _T_1619; // @[Counter.scala 35:22:@814.6]
  wire [5:0] _GEN_0; // @[Counter.scala 37:21:@816.6]
  wire  _T_2365; // @[BrCondTests.scala 32:32:@1187.4]
  wire  _T_2367; // @[BrCondTests.scala 33:32:@1188.4]
  wire  _T_2369; // @[BrCondTests.scala 34:32:@1189.4]
  wire  _T_2371; // @[BrCondTests.scala 35:32:@1190.4]
  wire  _T_2373; // @[BrCondTests.scala 36:32:@1191.4]
  wire  _T_2375; // @[BrCondTests.scala 37:32:@1192.4]
  wire  _GEN_4; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_5; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_6; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_7; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_8; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_9; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_10; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_11; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_12; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_13; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_14; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_15; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_16; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_17; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_18; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_19; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_20; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_21; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_22; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_23; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_24; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_25; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_26; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_27; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_28; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_29; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_30; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_31; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_32; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_33; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_34; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_35; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_36; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_37; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_38; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_39; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_40; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_41; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_42; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_43; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_44; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_45; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_46; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_47; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_48; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_49; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_50; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_51; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_52; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_53; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_54; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_55; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_56; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_57; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_58; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_59; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_60; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_61; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _T_2378; // @[BrCondTests.scala 37:16:@1193.4]
  wire  _GEN_64; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_65; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_66; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_67; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_68; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_69; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_70; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_71; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_72; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_73; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_74; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_75; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_76; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_77; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_78; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_79; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_80; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_81; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_82; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_83; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_84; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_85; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_86; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_87; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_88; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_89; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_90; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_91; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_92; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_93; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_94; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_95; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_96; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_97; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_98; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_99; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_100; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_101; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_102; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_103; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_104; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_105; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_106; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_107; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_108; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_109; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_110; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_111; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_112; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_113; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_114; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_115; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_116; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_117; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_118; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_119; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_120; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_121; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _T_2379; // @[BrCondTests.scala 36:16:@1194.4]
  wire  _GEN_123; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_124; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_125; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_126; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_127; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_128; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_129; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_130; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_131; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_132; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_133; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_134; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_135; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_136; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_137; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_138; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_139; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_140; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_141; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_142; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_143; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_144; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_145; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_146; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_147; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_148; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_149; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_150; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_151; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_152; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_153; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_154; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_155; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_156; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_157; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_158; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_159; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_160; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_161; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_162; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_163; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_164; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_165; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_166; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_167; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_168; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_169; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_170; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_171; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_172; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_173; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_174; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_175; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_176; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_177; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_178; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_179; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_180; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_181; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _T_2380; // @[BrCondTests.scala 35:16:@1195.4]
  wire  _GEN_183; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_184; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_185; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_186; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_187; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_188; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_189; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_190; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_191; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_192; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_193; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_194; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_195; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_196; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_197; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_198; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_199; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_200; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_201; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_202; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_203; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_204; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_205; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_206; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_207; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_208; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_209; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_210; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_211; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_212; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_213; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_214; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_215; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_216; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_217; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_218; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_219; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_220; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_221; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_222; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_223; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_224; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_225; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_226; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_227; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_228; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_229; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_230; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_231; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_232; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_233; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_234; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_235; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_236; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_237; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_238; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_239; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_240; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _GEN_241; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _T_2381; // @[BrCondTests.scala 34:16:@1196.4]
  wire  _T_2382; // @[BrCondTests.scala 33:16:@1197.4]
  wire  out; // @[BrCondTests.scala 32:16:@1198.4]
  wire [31:0] _GEN_363; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_364; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_365; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_366; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_367; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_368; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_369; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_370; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_371; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_372; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_373; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_374; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_375; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_376; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_377; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_378; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_379; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_380; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_381; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_382; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_383; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_384; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_385; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_386; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_387; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_388; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_389; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_390; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_391; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_392; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_393; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_394; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_395; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_396; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_397; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_398; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_399; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_400; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_401; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_402; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_403; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_404; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_405; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_406; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_407; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_408; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_409; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_410; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_411; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_412; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_413; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_414; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_415; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_416; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_417; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_418; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_419; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_420; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_421; // @[BrCondTests.scala 39:16:@1260.4]
  wire [31:0] _GEN_423; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_424; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_425; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_426; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_427; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_428; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_429; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_430; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_431; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_432; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_433; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_434; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_435; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_436; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_437; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_438; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_439; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_440; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_441; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_442; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_443; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_444; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_445; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_446; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_447; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_448; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_449; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_450; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_451; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_452; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_453; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_454; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_455; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_456; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_457; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_458; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_459; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_460; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_461; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_462; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_463; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_464; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_465; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_466; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_467; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_468; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_469; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_470; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_471; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_472; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_473; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_474; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_475; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_476; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_477; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_478; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_479; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_480; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_481; // @[BrCondTests.scala 41:14:@1323.4]
  wire [31:0] _GEN_483; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_484; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_485; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_486; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_487; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_488; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_489; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_490; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_491; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_492; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_493; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_494; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_495; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_496; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_497; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_498; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_499; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_500; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_501; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_502; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_503; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_504; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_505; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_506; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_507; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_508; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_509; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_510; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_511; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_512; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_513; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_514; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_515; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_516; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_517; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_518; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_519; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_520; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_521; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_522; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_523; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_524; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_525; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_526; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_527; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_528; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_529; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_530; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_531; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_532; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_533; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_534; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_535; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_536; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_537; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_538; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_539; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_540; // @[BrCondTests.scala 42:14:@1385.4]
  wire [31:0] _GEN_541; // @[BrCondTests.scala 42:14:@1385.4]
  wire  _T_2703; // @[BrCondTests.scala 44:20:@1388.6]
  wire  _T_2707; // @[BrCondTests.scala 45:23:@1398.4]
  wire  _T_2709; // @[BrCondTests.scala 45:9:@1400.4]
  wire  _T_2711; // @[BrCondTests.scala 45:9:@1401.4]
  BrCondArea dut ( // @[BrCondTests.scala 11:19:@804.4]
    .io_rs1(dut_io_rs1),
    .io_rs2(dut_io_rs2),
    .io_br_type(dut_io_br_type),
    .io_taken(dut_io_taken)
  );
  Control ctrl ( // @[BrCondTests.scala 12:20:@807.4]
    .io_inst(ctrl_io_inst),
    .io_br_type(ctrl_io_br_type)
  );
  assign done = value == 6'h3b; // @[Counter.scala 34:24:@812.6]
  assign _T_1618 = value + 6'h1; // @[Counter.scala 35:22:@813.6]
  assign _T_1619 = _T_1618[5:0]; // @[Counter.scala 35:22:@814.6]
  assign _GEN_0 = done ? 6'h0 : _T_1619; // @[Counter.scala 37:21:@816.6]
  assign _T_2365 = dut_io_br_type == 3'h3; // @[BrCondTests.scala 32:32:@1187.4]
  assign _T_2367 = dut_io_br_type == 3'h6; // @[BrCondTests.scala 33:32:@1188.4]
  assign _T_2369 = dut_io_br_type == 3'h2; // @[BrCondTests.scala 34:32:@1189.4]
  assign _T_2371 = dut_io_br_type == 3'h5; // @[BrCondTests.scala 35:32:@1190.4]
  assign _T_2373 = dut_io_br_type == 3'h1; // @[BrCondTests.scala 36:32:@1191.4]
  assign _T_2375 = dut_io_br_type == 3'h4; // @[BrCondTests.scala 37:32:@1192.4]
  assign _GEN_4 = 6'h2 == value ? 1'h0 : 1'h1; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_5 = 6'h3 == value ? 1'h0 : _GEN_4; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_6 = 6'h4 == value ? 1'h0 : _GEN_5; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_7 = 6'h5 == value ? 1'h0 : _GEN_6; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_8 = 6'h6 == value ? 1'h1 : _GEN_7; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_9 = 6'h7 == value ? 1'h1 : _GEN_8; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_10 = 6'h8 == value ? 1'h1 : _GEN_9; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_11 = 6'h9 == value ? 1'h1 : _GEN_10; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_12 = 6'ha == value ? 1'h1 : _GEN_11; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_13 = 6'hb == value ? 1'h1 : _GEN_12; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_14 = 6'hc == value ? 1'h0 : _GEN_13; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_15 = 6'hd == value ? 1'h0 : _GEN_14; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_16 = 6'he == value ? 1'h1 : _GEN_15; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_17 = 6'hf == value ? 1'h0 : _GEN_16; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_18 = 6'h10 == value ? 1'h1 : _GEN_17; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_19 = 6'h11 == value ? 1'h0 : _GEN_18; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_20 = 6'h12 == value ? 1'h1 : _GEN_19; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_21 = 6'h13 == value ? 1'h1 : _GEN_20; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_22 = 6'h14 == value ? 1'h0 : _GEN_21; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_23 = 6'h15 == value ? 1'h0 : _GEN_22; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_24 = 6'h16 == value ? 1'h1 : _GEN_23; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_25 = 6'h17 == value ? 1'h1 : _GEN_24; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_26 = 6'h18 == value ? 1'h0 : _GEN_25; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_27 = 6'h19 == value ? 1'h0 : _GEN_26; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_28 = 6'h1a == value ? 1'h0 : _GEN_27; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_29 = 6'h1b == value ? 1'h0 : _GEN_28; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_30 = 6'h1c == value ? 1'h1 : _GEN_29; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_31 = 6'h1d == value ? 1'h0 : _GEN_30; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_32 = 6'h1e == value ? 1'h1 : _GEN_31; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_33 = 6'h1f == value ? 1'h0 : _GEN_32; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_34 = 6'h20 == value ? 1'h1 : _GEN_33; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_35 = 6'h21 == value ? 1'h0 : _GEN_34; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_36 = 6'h22 == value ? 1'h0 : _GEN_35; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_37 = 6'h23 == value ? 1'h0 : _GEN_36; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_38 = 6'h24 == value ? 1'h0 : _GEN_37; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_39 = 6'h25 == value ? 1'h1 : _GEN_38; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_40 = 6'h26 == value ? 1'h1 : _GEN_39; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_41 = 6'h27 == value ? 1'h0 : _GEN_40; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_42 = 6'h28 == value ? 1'h1 : _GEN_41; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_43 = 6'h29 == value ? 1'h1 : _GEN_42; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_44 = 6'h2a == value ? 1'h0 : _GEN_43; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_45 = 6'h2b == value ? 1'h0 : _GEN_44; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_46 = 6'h2c == value ? 1'h1 : _GEN_45; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_47 = 6'h2d == value ? 1'h1 : _GEN_46; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_48 = 6'h2e == value ? 1'h1 : _GEN_47; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_49 = 6'h2f == value ? 1'h0 : _GEN_48; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_50 = 6'h30 == value ? 1'h0 : _GEN_49; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_51 = 6'h31 == value ? 1'h1 : _GEN_50; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_52 = 6'h32 == value ? 1'h0 : _GEN_51; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_53 = 6'h33 == value ? 1'h1 : _GEN_52; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_54 = 6'h34 == value ? 1'h0 : _GEN_53; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_55 = 6'h35 == value ? 1'h1 : _GEN_54; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_56 = 6'h36 == value ? 1'h0 : _GEN_55; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_57 = 6'h37 == value ? 1'h0 : _GEN_56; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_58 = 6'h38 == value ? 1'h0 : _GEN_57; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_59 = 6'h39 == value ? 1'h0 : _GEN_58; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_60 = 6'h3a == value ? 1'h0 : _GEN_59; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_61 = 6'h3b == value ? 1'h0 : _GEN_60; // @[BrCondTests.scala 37:16:@1193.4]
  assign _T_2378 = _T_2375 ? _GEN_61 : 1'h0; // @[BrCondTests.scala 37:16:@1193.4]
  assign _GEN_64 = 6'h2 == value; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_65 = 6'h3 == value ? 1'h1 : _GEN_64; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_66 = 6'h4 == value ? 1'h1 : _GEN_65; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_67 = 6'h5 == value ? 1'h1 : _GEN_66; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_68 = 6'h6 == value ? 1'h0 : _GEN_67; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_69 = 6'h7 == value ? 1'h0 : _GEN_68; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_70 = 6'h8 == value ? 1'h0 : _GEN_69; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_71 = 6'h9 == value ? 1'h0 : _GEN_70; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_72 = 6'ha == value ? 1'h0 : _GEN_71; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_73 = 6'hb == value ? 1'h0 : _GEN_72; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_74 = 6'hc == value ? 1'h1 : _GEN_73; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_75 = 6'hd == value ? 1'h1 : _GEN_74; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_76 = 6'he == value ? 1'h0 : _GEN_75; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_77 = 6'hf == value ? 1'h1 : _GEN_76; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_78 = 6'h10 == value ? 1'h0 : _GEN_77; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_79 = 6'h11 == value ? 1'h1 : _GEN_78; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_80 = 6'h12 == value ? 1'h0 : _GEN_79; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_81 = 6'h13 == value ? 1'h0 : _GEN_80; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_82 = 6'h14 == value ? 1'h1 : _GEN_81; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_83 = 6'h15 == value ? 1'h1 : _GEN_82; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_84 = 6'h16 == value ? 1'h0 : _GEN_83; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_85 = 6'h17 == value ? 1'h0 : _GEN_84; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_86 = 6'h18 == value ? 1'h1 : _GEN_85; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_87 = 6'h19 == value ? 1'h1 : _GEN_86; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_88 = 6'h1a == value ? 1'h1 : _GEN_87; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_89 = 6'h1b == value ? 1'h1 : _GEN_88; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_90 = 6'h1c == value ? 1'h0 : _GEN_89; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_91 = 6'h1d == value ? 1'h1 : _GEN_90; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_92 = 6'h1e == value ? 1'h0 : _GEN_91; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_93 = 6'h1f == value ? 1'h1 : _GEN_92; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_94 = 6'h20 == value ? 1'h0 : _GEN_93; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_95 = 6'h21 == value ? 1'h1 : _GEN_94; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_96 = 6'h22 == value ? 1'h1 : _GEN_95; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_97 = 6'h23 == value ? 1'h1 : _GEN_96; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_98 = 6'h24 == value ? 1'h1 : _GEN_97; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_99 = 6'h25 == value ? 1'h0 : _GEN_98; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_100 = 6'h26 == value ? 1'h0 : _GEN_99; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_101 = 6'h27 == value ? 1'h1 : _GEN_100; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_102 = 6'h28 == value ? 1'h0 : _GEN_101; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_103 = 6'h29 == value ? 1'h0 : _GEN_102; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_104 = 6'h2a == value ? 1'h1 : _GEN_103; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_105 = 6'h2b == value ? 1'h1 : _GEN_104; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_106 = 6'h2c == value ? 1'h0 : _GEN_105; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_107 = 6'h2d == value ? 1'h0 : _GEN_106; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_108 = 6'h2e == value ? 1'h0 : _GEN_107; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_109 = 6'h2f == value ? 1'h1 : _GEN_108; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_110 = 6'h30 == value ? 1'h1 : _GEN_109; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_111 = 6'h31 == value ? 1'h0 : _GEN_110; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_112 = 6'h32 == value ? 1'h1 : _GEN_111; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_113 = 6'h33 == value ? 1'h0 : _GEN_112; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_114 = 6'h34 == value ? 1'h1 : _GEN_113; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_115 = 6'h35 == value ? 1'h0 : _GEN_114; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_116 = 6'h36 == value ? 1'h1 : _GEN_115; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_117 = 6'h37 == value ? 1'h1 : _GEN_116; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_118 = 6'h38 == value ? 1'h1 : _GEN_117; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_119 = 6'h39 == value ? 1'h1 : _GEN_118; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_120 = 6'h3a == value ? 1'h1 : _GEN_119; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_121 = 6'h3b == value ? 1'h1 : _GEN_120; // @[BrCondTests.scala 36:16:@1194.4]
  assign _T_2379 = _T_2373 ? _GEN_121 : _T_2378; // @[BrCondTests.scala 36:16:@1194.4]
  assign _GEN_123 = 6'h1 == value ? 1'h0 : 1'h1; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_124 = 6'h2 == value ? 1'h0 : _GEN_123; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_125 = 6'h3 == value ? 1'h0 : _GEN_124; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_126 = 6'h4 == value ? 1'h0 : _GEN_125; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_127 = 6'h5 == value ? 1'h0 : _GEN_126; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_128 = 6'h6 == value ? 1'h1 : _GEN_127; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_129 = 6'h7 == value ? 1'h1 : _GEN_128; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_130 = 6'h8 == value ? 1'h0 : _GEN_129; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_131 = 6'h9 == value ? 1'h1 : _GEN_130; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_132 = 6'ha == value ? 1'h1 : _GEN_131; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_133 = 6'hb == value ? 1'h1 : _GEN_132; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_134 = 6'hc == value ? 1'h1 : _GEN_133; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_135 = 6'hd == value ? 1'h1 : _GEN_134; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_136 = 6'he == value ? 1'h1 : _GEN_135; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_137 = 6'hf == value ? 1'h1 : _GEN_136; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_138 = 6'h10 == value ? 1'h0 : _GEN_137; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_139 = 6'h11 == value ? 1'h1 : _GEN_138; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_140 = 6'h12 == value ? 1'h0 : _GEN_139; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_141 = 6'h13 == value ? 1'h0 : _GEN_140; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_142 = 6'h14 == value ? 1'h0 : _GEN_141; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_143 = 6'h15 == value ? 1'h1 : _GEN_142; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_144 = 6'h16 == value ? 1'h1 : _GEN_143; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_145 = 6'h17 == value ? 1'h0 : _GEN_144; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_146 = 6'h18 == value ? 1'h0 : _GEN_145; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_147 = 6'h19 == value ? 1'h0 : _GEN_146; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_148 = 6'h1a == value ? 1'h0 : _GEN_147; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_149 = 6'h1b == value ? 1'h1 : _GEN_148; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_150 = 6'h1c == value ? 1'h1 : _GEN_149; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_151 = 6'h1d == value ? 1'h1 : _GEN_150; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_152 = 6'h1e == value ? 1'h0 : _GEN_151; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_153 = 6'h1f == value ? 1'h1 : _GEN_152; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_154 = 6'h20 == value ? 1'h1 : _GEN_153; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_155 = 6'h21 == value ? 1'h0 : _GEN_154; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_156 = 6'h22 == value ? 1'h0 : _GEN_155; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_157 = 6'h23 == value ? 1'h0 : _GEN_156; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_158 = 6'h24 == value ? 1'h0 : _GEN_157; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_159 = 6'h25 == value ? 1'h1 : _GEN_158; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_160 = 6'h26 == value ? 1'h0 : _GEN_159; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_161 = 6'h27 == value ? 1'h1 : _GEN_160; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_162 = 6'h28 == value ? 1'h1 : _GEN_161; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_163 = 6'h29 == value ? 1'h0 : _GEN_162; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_164 = 6'h2a == value ? 1'h0 : _GEN_163; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_165 = 6'h2b == value ? 1'h1 : _GEN_164; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_166 = 6'h2c == value ? 1'h1 : _GEN_165; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_167 = 6'h2d == value ? 1'h1 : _GEN_166; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_168 = 6'h2e == value ? 1'h1 : _GEN_167; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_169 = 6'h2f == value ? 1'h0 : _GEN_168; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_170 = 6'h30 == value ? 1'h0 : _GEN_169; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_171 = 6'h31 == value ? 1'h1 : _GEN_170; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_172 = 6'h32 == value ? 1'h0 : _GEN_171; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_173 = 6'h33 == value ? 1'h1 : _GEN_172; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_174 = 6'h34 == value ? 1'h1 : _GEN_173; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_175 = 6'h35 == value ? 1'h0 : _GEN_174; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_176 = 6'h36 == value ? 1'h1 : _GEN_175; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_177 = 6'h37 == value ? 1'h1 : _GEN_176; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_178 = 6'h38 == value ? 1'h1 : _GEN_177; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_179 = 6'h39 == value ? 1'h1 : _GEN_178; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_180 = 6'h3a == value ? 1'h0 : _GEN_179; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_181 = 6'h3b == value ? 1'h0 : _GEN_180; // @[BrCondTests.scala 35:16:@1195.4]
  assign _T_2380 = _T_2371 ? _GEN_181 : _T_2379; // @[BrCondTests.scala 35:16:@1195.4]
  assign _GEN_183 = 6'h1 == value; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_184 = 6'h2 == value ? 1'h1 : _GEN_183; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_185 = 6'h3 == value ? 1'h1 : _GEN_184; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_186 = 6'h4 == value ? 1'h1 : _GEN_185; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_187 = 6'h5 == value ? 1'h1 : _GEN_186; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_188 = 6'h6 == value ? 1'h0 : _GEN_187; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_189 = 6'h7 == value ? 1'h0 : _GEN_188; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_190 = 6'h8 == value ? 1'h1 : _GEN_189; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_191 = 6'h9 == value ? 1'h0 : _GEN_190; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_192 = 6'ha == value ? 1'h0 : _GEN_191; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_193 = 6'hb == value ? 1'h0 : _GEN_192; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_194 = 6'hc == value ? 1'h0 : _GEN_193; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_195 = 6'hd == value ? 1'h0 : _GEN_194; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_196 = 6'he == value ? 1'h0 : _GEN_195; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_197 = 6'hf == value ? 1'h0 : _GEN_196; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_198 = 6'h10 == value ? 1'h1 : _GEN_197; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_199 = 6'h11 == value ? 1'h0 : _GEN_198; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_200 = 6'h12 == value ? 1'h1 : _GEN_199; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_201 = 6'h13 == value ? 1'h1 : _GEN_200; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_202 = 6'h14 == value ? 1'h1 : _GEN_201; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_203 = 6'h15 == value ? 1'h0 : _GEN_202; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_204 = 6'h16 == value ? 1'h0 : _GEN_203; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_205 = 6'h17 == value ? 1'h1 : _GEN_204; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_206 = 6'h18 == value ? 1'h1 : _GEN_205; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_207 = 6'h19 == value ? 1'h1 : _GEN_206; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_208 = 6'h1a == value ? 1'h1 : _GEN_207; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_209 = 6'h1b == value ? 1'h0 : _GEN_208; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_210 = 6'h1c == value ? 1'h0 : _GEN_209; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_211 = 6'h1d == value ? 1'h0 : _GEN_210; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_212 = 6'h1e == value ? 1'h1 : _GEN_211; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_213 = 6'h1f == value ? 1'h0 : _GEN_212; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_214 = 6'h20 == value ? 1'h0 : _GEN_213; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_215 = 6'h21 == value ? 1'h1 : _GEN_214; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_216 = 6'h22 == value ? 1'h1 : _GEN_215; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_217 = 6'h23 == value ? 1'h1 : _GEN_216; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_218 = 6'h24 == value ? 1'h1 : _GEN_217; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_219 = 6'h25 == value ? 1'h0 : _GEN_218; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_220 = 6'h26 == value ? 1'h1 : _GEN_219; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_221 = 6'h27 == value ? 1'h0 : _GEN_220; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_222 = 6'h28 == value ? 1'h0 : _GEN_221; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_223 = 6'h29 == value ? 1'h1 : _GEN_222; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_224 = 6'h2a == value ? 1'h1 : _GEN_223; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_225 = 6'h2b == value ? 1'h0 : _GEN_224; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_226 = 6'h2c == value ? 1'h0 : _GEN_225; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_227 = 6'h2d == value ? 1'h0 : _GEN_226; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_228 = 6'h2e == value ? 1'h0 : _GEN_227; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_229 = 6'h2f == value ? 1'h1 : _GEN_228; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_230 = 6'h30 == value ? 1'h1 : _GEN_229; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_231 = 6'h31 == value ? 1'h0 : _GEN_230; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_232 = 6'h32 == value ? 1'h1 : _GEN_231; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_233 = 6'h33 == value ? 1'h0 : _GEN_232; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_234 = 6'h34 == value ? 1'h0 : _GEN_233; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_235 = 6'h35 == value ? 1'h1 : _GEN_234; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_236 = 6'h36 == value ? 1'h0 : _GEN_235; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_237 = 6'h37 == value ? 1'h0 : _GEN_236; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_238 = 6'h38 == value ? 1'h0 : _GEN_237; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_239 = 6'h39 == value ? 1'h0 : _GEN_238; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_240 = 6'h3a == value ? 1'h1 : _GEN_239; // @[BrCondTests.scala 34:16:@1196.4]
  assign _GEN_241 = 6'h3b == value ? 1'h1 : _GEN_240; // @[BrCondTests.scala 34:16:@1196.4]
  assign _T_2381 = _T_2369 ? _GEN_241 : _T_2380; // @[BrCondTests.scala 34:16:@1196.4]
  assign _T_2382 = _T_2367 ? 1'h1 : _T_2381; // @[BrCondTests.scala 33:16:@1197.4]
  assign out = _T_2365 ? 1'h0 : _T_2382; // @[BrCondTests.scala 32:16:@1198.4]
  assign _GEN_363 = 6'h1 == value ? 32'h1063 : 32'h63; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_364 = 6'h2 == value ? 32'h4063 : _GEN_363; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_365 = 6'h3 == value ? 32'h5063 : _GEN_364; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_366 = 6'h4 == value ? 32'h6063 : _GEN_365; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_367 = 6'h5 == value ? 32'h7063 : _GEN_366; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_368 = 6'h6 == value ? 32'h63 : _GEN_367; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_369 = 6'h7 == value ? 32'h1063 : _GEN_368; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_370 = 6'h8 == value ? 32'h4063 : _GEN_369; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_371 = 6'h9 == value ? 32'h5063 : _GEN_370; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_372 = 6'ha == value ? 32'h6063 : _GEN_371; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_373 = 6'hb == value ? 32'h7063 : _GEN_372; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_374 = 6'hc == value ? 32'h63 : _GEN_373; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_375 = 6'hd == value ? 32'h1063 : _GEN_374; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_376 = 6'he == value ? 32'h4063 : _GEN_375; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_377 = 6'hf == value ? 32'h5063 : _GEN_376; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_378 = 6'h10 == value ? 32'h6063 : _GEN_377; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_379 = 6'h11 == value ? 32'h7063 : _GEN_378; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_380 = 6'h12 == value ? 32'h63 : _GEN_379; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_381 = 6'h13 == value ? 32'h1063 : _GEN_380; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_382 = 6'h14 == value ? 32'h4063 : _GEN_381; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_383 = 6'h15 == value ? 32'h5063 : _GEN_382; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_384 = 6'h16 == value ? 32'h6063 : _GEN_383; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_385 = 6'h17 == value ? 32'h7063 : _GEN_384; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_386 = 6'h18 == value ? 32'h63 : _GEN_385; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_387 = 6'h19 == value ? 32'h1063 : _GEN_386; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_388 = 6'h1a == value ? 32'h4063 : _GEN_387; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_389 = 6'h1b == value ? 32'h5063 : _GEN_388; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_390 = 6'h1c == value ? 32'h6063 : _GEN_389; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_391 = 6'h1d == value ? 32'h7063 : _GEN_390; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_392 = 6'h1e == value ? 32'h63 : _GEN_391; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_393 = 6'h1f == value ? 32'h1063 : _GEN_392; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_394 = 6'h20 == value ? 32'h4063 : _GEN_393; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_395 = 6'h21 == value ? 32'h5063 : _GEN_394; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_396 = 6'h22 == value ? 32'h6063 : _GEN_395; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_397 = 6'h23 == value ? 32'h7063 : _GEN_396; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_398 = 6'h24 == value ? 32'h63 : _GEN_397; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_399 = 6'h25 == value ? 32'h1063 : _GEN_398; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_400 = 6'h26 == value ? 32'h4063 : _GEN_399; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_401 = 6'h27 == value ? 32'h5063 : _GEN_400; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_402 = 6'h28 == value ? 32'h6063 : _GEN_401; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_403 = 6'h29 == value ? 32'h7063 : _GEN_402; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_404 = 6'h2a == value ? 32'h63 : _GEN_403; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_405 = 6'h2b == value ? 32'h1063 : _GEN_404; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_406 = 6'h2c == value ? 32'h4063 : _GEN_405; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_407 = 6'h2d == value ? 32'h5063 : _GEN_406; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_408 = 6'h2e == value ? 32'h6063 : _GEN_407; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_409 = 6'h2f == value ? 32'h7063 : _GEN_408; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_410 = 6'h30 == value ? 32'h63 : _GEN_409; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_411 = 6'h31 == value ? 32'h1063 : _GEN_410; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_412 = 6'h32 == value ? 32'h4063 : _GEN_411; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_413 = 6'h33 == value ? 32'h5063 : _GEN_412; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_414 = 6'h34 == value ? 32'h6063 : _GEN_413; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_415 = 6'h35 == value ? 32'h7063 : _GEN_414; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_416 = 6'h36 == value ? 32'h63 : _GEN_415; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_417 = 6'h37 == value ? 32'h1063 : _GEN_416; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_418 = 6'h38 == value ? 32'h4063 : _GEN_417; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_419 = 6'h39 == value ? 32'h5063 : _GEN_418; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_420 = 6'h3a == value ? 32'h6063 : _GEN_419; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_421 = 6'h3b == value ? 32'h7063 : _GEN_420; // @[BrCondTests.scala 39:16:@1260.4]
  assign _GEN_423 = 6'h1 == value ? 32'heedc498d : 32'h1b5c55a; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_424 = 6'h2 == value ? 32'h86f8a91d : _GEN_423; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_425 = 6'h3 == value ? 32'h8fda0b0e : _GEN_424; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_426 = 6'h4 == value ? 32'h1a727694 : _GEN_425; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_427 = 6'h5 == value ? 32'h8ab69259 : _GEN_426; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_428 = 6'h6 == value ? 32'h5e476af2 : _GEN_427; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_429 = 6'h7 == value ? 32'hf81e7dc2 : _GEN_428; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_430 = 6'h8 == value ? 32'hc15dc176 : _GEN_429; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_431 = 6'h9 == value ? 32'h6b8383ff : _GEN_430; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_432 = 6'ha == value ? 32'h3114f9d7 : _GEN_431; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_433 = 6'hb == value ? 32'h3c3794cc : _GEN_432; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_434 = 6'hc == value ? 32'hf5dbfcb : _GEN_433; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_435 = 6'hd == value ? 32'h608fd458 : _GEN_434; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_436 = 6'he == value ? 32'h6c9f5cc6 : _GEN_435; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_437 = 6'hf == value ? 32'h392bd9d5 : _GEN_436; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_438 = 6'h10 == value ? 32'h8d309823 : _GEN_437; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_439 = 6'h11 == value ? 32'h491c13de : _GEN_438; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_440 = 6'h12 == value ? 32'he0797750 : _GEN_439; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_441 = 6'h13 == value ? 32'hef68d993 : _GEN_440; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_442 = 6'h14 == value ? 32'h11f8bec3 : _GEN_441; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_443 = 6'h15 == value ? 32'h515f8d94 : _GEN_442; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_444 = 6'h16 == value ? 32'h6c1b35ae : _GEN_443; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_445 = 6'h17 == value ? 32'heb2fe04b : _GEN_444; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_446 = 6'h18 == value ? 32'h2c97d1db : _GEN_445; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_447 = 6'h19 == value ? 32'h87fec123 : _GEN_446; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_448 = 6'h1a == value ? 32'he53fe615 : _GEN_447; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_449 = 6'h1b == value ? 32'h50737a97 : _GEN_448; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_450 = 6'h1c == value ? 32'hdf5e84fe : _GEN_449; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_451 = 6'h1d == value ? 32'h7c6cdb45 : _GEN_450; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_452 = 6'h1e == value ? 32'hcdc0534e : _GEN_451; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_453 = 6'h1f == value ? 32'h1505be69 : _GEN_452; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_454 = 6'h20 == value ? 32'hc30b4fce : _GEN_453; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_455 = 6'h21 == value ? 32'h1c41d066 : _GEN_454; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_456 = 6'h22 == value ? 32'hb45b7485 : _GEN_455; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_457 = 6'h23 == value ? 32'h7373a04f : _GEN_456; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_458 = 6'h24 == value ? 32'h8f78d3f6 : _GEN_457; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_459 = 6'h25 == value ? 32'h2a04fd88 : _GEN_458; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_460 = 6'h26 == value ? 32'hdfb9c660 : _GEN_459; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_461 = 6'h27 == value ? 32'h33e9d8f8 : _GEN_460; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_462 = 6'h28 == value ? 32'hd8f82e5d : _GEN_461; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_463 = 6'h29 == value ? 32'hf5867366 : _GEN_462; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_464 = 6'h2a == value ? 32'h8324a153 : _GEN_463; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_465 = 6'h2b == value ? 32'h43441ef6 : _GEN_464; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_466 = 6'h2c == value ? 32'h4862a797 : _GEN_465; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_467 = 6'h2d == value ? 32'h62df4fdc : _GEN_466; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_468 = 6'h2e == value ? 32'h2a2c2132 : _GEN_467; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_469 = 6'h2f == value ? 32'h6b2fb8c4 : _GEN_468; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_470 = 6'h30 == value ? 32'h24b1779f : _GEN_469; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_471 = 6'h31 == value ? 32'h5bd3c985 : _GEN_470; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_472 = 6'h32 == value ? 32'h90b7207 : _GEN_471; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_473 = 6'h33 == value ? 32'h5556ab0b : _GEN_472; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_474 = 6'h34 == value ? 32'h16a190c3 : _GEN_473; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_475 = 6'h35 == value ? 32'hf5d7d1a5 : _GEN_474; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_476 = 6'h36 == value ? 32'h4c449625 : _GEN_475; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_477 = 6'h37 == value ? 32'h57190720 : _GEN_476; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_478 = 6'h38 == value ? 32'h3cd4a5df : _GEN_477; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_479 = 6'h39 == value ? 32'h7fa17049 : _GEN_478; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_480 = 6'h3a == value ? 32'h87e9f97d : _GEN_479; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_481 = 6'h3b == value ? 32'h97ae1dd1 : _GEN_480; // @[BrCondTests.scala 41:14:@1323.4]
  assign _GEN_483 = 6'h1 == value ? 32'h4a423ead : 32'h3fdfcd; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_484 = 6'h2 == value ? 32'hc79d662f : _GEN_483; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_485 = 6'h3 == value ? 32'hbfdf9a61 : _GEN_484; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_486 = 6'h4 == value ? 32'h60cbf61b : _GEN_485; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_487 = 6'h5 == value ? 32'hfd73a3dd : _GEN_486; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_488 = 6'h6 == value ? 32'h10b12e64 : _GEN_487; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_489 = 6'h7 == value ? 32'h952cc9d0 : _GEN_488; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_490 = 6'h8 == value ? 32'h60119efe : _GEN_489; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_491 = 6'h9 == value ? 32'h2357b79e : _GEN_490; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_492 = 6'ha == value ? 32'h11519f5a : _GEN_491; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_493 = 6'hb == value ? 32'h3a44925e : _GEN_492; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_494 = 6'hc == value ? 32'haf588a87 : _GEN_493; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_495 = 6'hd == value ? 32'hffaaef8d : _GEN_494; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_496 = 6'he == value ? 32'h376a11bf : _GEN_495; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_497 = 6'hf == value ? 32'ha0a8df52 : _GEN_496; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_498 = 6'h10 == value ? 32'h35ae5d14 : _GEN_497; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_499 = 6'h11 == value ? 32'hc780fa89 : _GEN_498; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_500 = 6'h12 == value ? 32'h115a2b43 : _GEN_499; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_501 = 6'h13 == value ? 32'h5b3684f7 : _GEN_500; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_502 = 6'h14 == value ? 32'h764e5d08 : _GEN_501; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_503 = 6'h15 == value ? 32'h9b696e4e : _GEN_502; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_504 = 6'h16 == value ? 32'hec52568 : _GEN_503; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_505 = 6'h17 == value ? 32'h1378e0e7 : _GEN_504; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_506 = 6'h18 == value ? 32'h5de9c7be : _GEN_505; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_507 = 6'h19 == value ? 32'hd47f2b62 : _GEN_506; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_508 = 6'h1a == value ? 32'hf20e2d9c : _GEN_507; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_509 = 6'h1b == value ? 32'h8460ba8b : _GEN_508; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_510 = 6'h1c == value ? 32'hc1ec01ba : _GEN_509; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_511 = 6'h1d == value ? 32'hffaf9b33 : _GEN_510; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_512 = 6'h1e == value ? 32'h50b23288 : _GEN_511; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_513 = 6'h1f == value ? 32'hf06a27e1 : _GEN_512; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_514 = 6'h20 == value ? 32'h96d51621 : _GEN_513; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_515 = 6'h21 == value ? 32'h67b52c81 : _GEN_514; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_516 = 6'h22 == value ? 32'hc2e0b2aa : _GEN_515; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_517 = 6'h23 == value ? 32'h77b57a80 : _GEN_516; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_518 = 6'h24 == value ? 32'hf578396b : _GEN_517; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_519 = 6'h25 == value ? 32'h1012b1f9 : _GEN_518; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_520 = 6'h26 == value ? 32'heba6021 : _GEN_519; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_521 = 6'h27 == value ? 32'ha85378d9 : _GEN_520; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_522 = 6'h28 == value ? 32'hc9934356 : _GEN_521; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_523 = 6'h29 == value ? 32'h28138722 : _GEN_522; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_524 = 6'h2a == value ? 32'hfab5adc7 : _GEN_523; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_525 = 6'h2b == value ? 32'hd04567be : _GEN_524; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_526 = 6'h2c == value ? 32'h20f541d : _GEN_525; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_527 = 6'h2d == value ? 32'heae9f7c : _GEN_526; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_528 = 6'h2e == value ? 32'h22169984 : _GEN_527; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_529 = 6'h2f == value ? 32'h71b5a828 : _GEN_528; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_530 = 6'h30 == value ? 32'h538a18e9 : _GEN_529; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_531 = 6'h31 == value ? 32'h2d68e3e6 : _GEN_530; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_532 = 6'h32 == value ? 32'h576847e1 : _GEN_531; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_533 = 6'h33 == value ? 32'h36f5ed34 : _GEN_532; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_534 = 6'h34 == value ? 32'hc3ca6388 : _GEN_533; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_535 = 6'h35 == value ? 32'hb358240 : _GEN_534; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_536 = 6'h36 == value ? 32'hd8bc44db : _GEN_535; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_537 = 6'h37 == value ? 32'ha11c4e6f : _GEN_536; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_538 = 6'h38 == value ? 32'hefba095c : _GEN_537; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_539 = 6'h39 == value ? 32'hb7191350 : _GEN_538; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_540 = 6'h3a == value ? 32'hf15c7df9 : _GEN_539; // @[BrCondTests.scala 42:14:@1385.4]
  assign _GEN_541 = 6'h3b == value ? 32'ha9e8ba52 : _GEN_540; // @[BrCondTests.scala 42:14:@1385.4]
  assign _T_2703 = reset == 1'h0; // @[BrCondTests.scala 44:20:@1388.6]
  assign _T_2707 = dut_io_taken == out; // @[BrCondTests.scala 45:23:@1398.4]
  assign _T_2709 = _T_2707 | reset; // @[BrCondTests.scala 45:9:@1400.4]
  assign _T_2711 = _T_2709 == 1'h0; // @[BrCondTests.scala 45:9:@1401.4]
  assign dut_io_rs1 = _GEN_481;
  assign dut_io_rs2 = _GEN_541;
  assign dut_io_br_type = ctrl_io_br_type;
  assign ctrl_io_inst = _GEN_421;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  value = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      value <= 6'h0;
    end else begin
      if (done) begin
        value <= 6'h0;
      end else begin
        value <= _T_1619;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (done & _T_2703) begin
          $finish; // @[BrCondTests.scala 44:20:@1390.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (done & _T_2703) begin
          $finish; // @[BrCondTests.scala 44:28:@1395.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2711) begin
          $fwrite(32'h80000002,"Assertion failed\n    at BrCondTests.scala:45 assert(dut.io.taken === out)\n"); // @[BrCondTests.scala 45:9:@1403.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2711) begin
          $fatal; // @[BrCondTests.scala 45:9:@1404.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2703) begin
          $fwrite(32'h80000002,"Counter: %d, BrType: 0x%h, rs1: 0x%h, rs2: 0x%h, Taken: %d ?= %d\n",value,dut_io_br_type,dut_io_rs1,dut_io_rs2,dut_io_taken,out); // @[BrCondTests.scala 46:9:@1409.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
