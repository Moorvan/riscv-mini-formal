module ALUArea( // @[:@3.2]
  input  [31:0] io_A, // @[:@6.4]
  input  [31:0] io_B, // @[:@6.4]
  input  [3:0]  io_alu_op, // @[:@6.4]
  output [31:0] io_out, // @[:@6.4]
  output [31:0] io_sum // @[:@6.4]
);
  wire  _T_15; // @[ALU.scala 59:33:@8.4]
  wire [32:0] _T_17; // @[ALU.scala 59:38:@9.4]
  wire [32:0] _T_18; // @[ALU.scala 59:38:@10.4]
  wire [31:0] _T_19; // @[ALU.scala 59:38:@11.4]
  wire [31:0] _T_20; // @[ALU.scala 59:23:@12.4]
  wire [32:0] _T_21; // @[ALU.scala 59:18:@13.4]
  wire [31:0] sum; // @[ALU.scala 59:18:@14.4]
  wire  _T_22; // @[ALU.scala 60:21:@15.4]
  wire  _T_23; // @[ALU.scala 60:38:@16.4]
  wire  _T_24; // @[ALU.scala 60:30:@17.4]
  wire  _T_25; // @[ALU.scala 60:51:@18.4]
  wire  _T_26; // @[ALU.scala 61:26:@19.4]
  wire  _T_29; // @[ALU.scala 61:16:@22.4]
  wire  cmp; // @[ALU.scala 60:16:@23.4]
  wire [4:0] shamt; // @[ALU.scala 62:20:@24.4]
  wire  _T_30; // @[ALU.scala 63:29:@25.4]
  wire [15:0] _T_35; // @[Bitwise.scala 103:21:@28.4]
  wire [31:0] _T_36; // @[Bitwise.scala 103:31:@29.4]
  wire [15:0] _T_37; // @[Bitwise.scala 103:46:@30.4]
  wire [31:0] _GEN_0; // @[Bitwise.scala 103:65:@31.4]
  wire [31:0] _T_38; // @[Bitwise.scala 103:65:@31.4]
  wire [31:0] _T_40; // @[Bitwise.scala 103:75:@33.4]
  wire [31:0] _T_41; // @[Bitwise.scala 103:39:@34.4]
  wire [23:0] _T_45; // @[Bitwise.scala 103:21:@38.4]
  wire [31:0] _GEN_1; // @[Bitwise.scala 103:31:@39.4]
  wire [31:0] _T_46; // @[Bitwise.scala 103:31:@39.4]
  wire [23:0] _T_47; // @[Bitwise.scala 103:46:@40.4]
  wire [31:0] _GEN_2; // @[Bitwise.scala 103:65:@41.4]
  wire [31:0] _T_48; // @[Bitwise.scala 103:65:@41.4]
  wire [31:0] _T_50; // @[Bitwise.scala 103:75:@43.4]
  wire [31:0] _T_51; // @[Bitwise.scala 103:39:@44.4]
  wire [27:0] _T_55; // @[Bitwise.scala 103:21:@48.4]
  wire [31:0] _GEN_3; // @[Bitwise.scala 103:31:@49.4]
  wire [31:0] _T_56; // @[Bitwise.scala 103:31:@49.4]
  wire [27:0] _T_57; // @[Bitwise.scala 103:46:@50.4]
  wire [31:0] _GEN_4; // @[Bitwise.scala 103:65:@51.4]
  wire [31:0] _T_58; // @[Bitwise.scala 103:65:@51.4]
  wire [31:0] _T_60; // @[Bitwise.scala 103:75:@53.4]
  wire [31:0] _T_61; // @[Bitwise.scala 103:39:@54.4]
  wire [29:0] _T_65; // @[Bitwise.scala 103:21:@58.4]
  wire [31:0] _GEN_5; // @[Bitwise.scala 103:31:@59.4]
  wire [31:0] _T_66; // @[Bitwise.scala 103:31:@59.4]
  wire [29:0] _T_67; // @[Bitwise.scala 103:46:@60.4]
  wire [31:0] _GEN_6; // @[Bitwise.scala 103:65:@61.4]
  wire [31:0] _T_68; // @[Bitwise.scala 103:65:@61.4]
  wire [31:0] _T_70; // @[Bitwise.scala 103:75:@63.4]
  wire [31:0] _T_71; // @[Bitwise.scala 103:39:@64.4]
  wire [30:0] _T_75; // @[Bitwise.scala 103:21:@68.4]
  wire [31:0] _GEN_7; // @[Bitwise.scala 103:31:@69.4]
  wire [31:0] _T_76; // @[Bitwise.scala 103:31:@69.4]
  wire [30:0] _T_77; // @[Bitwise.scala 103:46:@70.4]
  wire [31:0] _GEN_8; // @[Bitwise.scala 103:65:@71.4]
  wire [31:0] _T_78; // @[Bitwise.scala 103:65:@71.4]
  wire [31:0] _T_80; // @[Bitwise.scala 103:75:@73.4]
  wire [31:0] _T_81; // @[Bitwise.scala 103:39:@74.4]
  wire [31:0] shin; // @[ALU.scala 63:19:@75.4]
  wire  _T_83; // @[ALU.scala 64:41:@77.4]
  wire  _T_84; // @[ALU.scala 64:34:@78.4]
  wire [32:0] _T_85; // @[Cat.scala 30:58:@79.4]
  wire [32:0] _T_86; // @[ALU.scala 64:57:@80.4]
  wire [32:0] _T_87; // @[ALU.scala 64:64:@81.4]
  wire [31:0] shiftr; // @[ALU.scala 64:73:@82.4]
  wire [15:0] _T_92; // @[Bitwise.scala 103:21:@85.4]
  wire [31:0] _T_93; // @[Bitwise.scala 103:31:@86.4]
  wire [15:0] _T_94; // @[Bitwise.scala 103:46:@87.4]
  wire [31:0] _GEN_9; // @[Bitwise.scala 103:65:@88.4]
  wire [31:0] _T_95; // @[Bitwise.scala 103:65:@88.4]
  wire [31:0] _T_97; // @[Bitwise.scala 103:75:@90.4]
  wire [31:0] _T_98; // @[Bitwise.scala 103:39:@91.4]
  wire [23:0] _T_102; // @[Bitwise.scala 103:21:@95.4]
  wire [31:0] _GEN_10; // @[Bitwise.scala 103:31:@96.4]
  wire [31:0] _T_103; // @[Bitwise.scala 103:31:@96.4]
  wire [23:0] _T_104; // @[Bitwise.scala 103:46:@97.4]
  wire [31:0] _GEN_11; // @[Bitwise.scala 103:65:@98.4]
  wire [31:0] _T_105; // @[Bitwise.scala 103:65:@98.4]
  wire [31:0] _T_107; // @[Bitwise.scala 103:75:@100.4]
  wire [31:0] _T_108; // @[Bitwise.scala 103:39:@101.4]
  wire [27:0] _T_112; // @[Bitwise.scala 103:21:@105.4]
  wire [31:0] _GEN_12; // @[Bitwise.scala 103:31:@106.4]
  wire [31:0] _T_113; // @[Bitwise.scala 103:31:@106.4]
  wire [27:0] _T_114; // @[Bitwise.scala 103:46:@107.4]
  wire [31:0] _GEN_13; // @[Bitwise.scala 103:65:@108.4]
  wire [31:0] _T_115; // @[Bitwise.scala 103:65:@108.4]
  wire [31:0] _T_117; // @[Bitwise.scala 103:75:@110.4]
  wire [31:0] _T_118; // @[Bitwise.scala 103:39:@111.4]
  wire [29:0] _T_122; // @[Bitwise.scala 103:21:@115.4]
  wire [31:0] _GEN_14; // @[Bitwise.scala 103:31:@116.4]
  wire [31:0] _T_123; // @[Bitwise.scala 103:31:@116.4]
  wire [29:0] _T_124; // @[Bitwise.scala 103:46:@117.4]
  wire [31:0] _GEN_15; // @[Bitwise.scala 103:65:@118.4]
  wire [31:0] _T_125; // @[Bitwise.scala 103:65:@118.4]
  wire [31:0] _T_127; // @[Bitwise.scala 103:75:@120.4]
  wire [31:0] _T_128; // @[Bitwise.scala 103:39:@121.4]
  wire [30:0] _T_132; // @[Bitwise.scala 103:21:@125.4]
  wire [31:0] _GEN_16; // @[Bitwise.scala 103:31:@126.4]
  wire [31:0] _T_133; // @[Bitwise.scala 103:31:@126.4]
  wire [30:0] _T_134; // @[Bitwise.scala 103:46:@127.4]
  wire [31:0] _GEN_17; // @[Bitwise.scala 103:65:@128.4]
  wire [31:0] _T_135; // @[Bitwise.scala 103:65:@128.4]
  wire [31:0] _T_137; // @[Bitwise.scala 103:75:@130.4]
  wire [31:0] shiftl; // @[Bitwise.scala 103:39:@131.4]
  wire  _T_151; // @[ALU.scala 68:19:@132.4]
  wire  _T_152; // @[ALU.scala 68:44:@133.4]
  wire  _T_153; // @[ALU.scala 68:31:@134.4]
  wire  _T_154; // @[ALU.scala 69:19:@135.4]
  wire  _T_155; // @[ALU.scala 69:44:@136.4]
  wire  _T_156; // @[ALU.scala 69:31:@137.4]
  wire  _T_157; // @[ALU.scala 70:19:@138.4]
  wire  _T_158; // @[ALU.scala 70:44:@139.4]
  wire  _T_159; // @[ALU.scala 70:31:@140.4]
  wire  _T_160; // @[ALU.scala 71:19:@141.4]
  wire  _T_161; // @[ALU.scala 72:19:@142.4]
  wire [31:0] _T_162; // @[ALU.scala 72:38:@143.4]
  wire  _T_163; // @[ALU.scala 73:19:@144.4]
  wire [31:0] _T_164; // @[ALU.scala 73:38:@145.4]
  wire  _T_165; // @[ALU.scala 74:19:@146.4]
  wire [31:0] _T_166; // @[ALU.scala 74:38:@147.4]
  wire  _T_167; // @[ALU.scala 75:19:@148.4]
  wire [31:0] _T_168; // @[ALU.scala 75:8:@149.4]
  wire [31:0] _T_169; // @[ALU.scala 74:8:@150.4]
  wire [31:0] _T_170; // @[ALU.scala 73:8:@151.4]
  wire [31:0] _T_171; // @[ALU.scala 72:8:@152.4]
  wire [31:0] _T_172; // @[ALU.scala 71:8:@153.4]
  wire [31:0] _T_173; // @[ALU.scala 70:8:@154.4]
  wire [31:0] _T_174; // @[ALU.scala 69:8:@155.4]
  wire [31:0] out; // @[ALU.scala 68:8:@156.4]
  assign _T_15 = io_alu_op[0]; // @[ALU.scala 59:33:@8.4]
  assign _T_17 = 32'h0 - io_B; // @[ALU.scala 59:38:@9.4]
  assign _T_18 = $unsigned(_T_17); // @[ALU.scala 59:38:@10.4]
  assign _T_19 = _T_18[31:0]; // @[ALU.scala 59:38:@11.4]
  assign _T_20 = _T_15 ? _T_19 : io_B; // @[ALU.scala 59:23:@12.4]
  assign _T_21 = io_A + _T_20; // @[ALU.scala 59:18:@13.4]
  assign sum = _T_21[31:0]; // @[ALU.scala 59:18:@14.4]
  assign _T_22 = io_A[31]; // @[ALU.scala 60:21:@15.4]
  assign _T_23 = io_B[31]; // @[ALU.scala 60:38:@16.4]
  assign _T_24 = _T_22 == _T_23; // @[ALU.scala 60:30:@17.4]
  assign _T_25 = sum[31]; // @[ALU.scala 60:51:@18.4]
  assign _T_26 = io_alu_op[1]; // @[ALU.scala 61:26:@19.4]
  assign _T_29 = _T_26 ? _T_23 : _T_22; // @[ALU.scala 61:16:@22.4]
  assign cmp = _T_24 ? _T_25 : _T_29; // @[ALU.scala 60:16:@23.4]
  assign shamt = io_B[4:0]; // @[ALU.scala 62:20:@24.4]
  assign _T_30 = io_alu_op[3]; // @[ALU.scala 63:29:@25.4]
  assign _T_35 = io_A[31:16]; // @[Bitwise.scala 103:21:@28.4]
  assign _T_36 = {{16'd0}, _T_35}; // @[Bitwise.scala 103:31:@29.4]
  assign _T_37 = io_A[15:0]; // @[Bitwise.scala 103:46:@30.4]
  assign _GEN_0 = {{16'd0}, _T_37}; // @[Bitwise.scala 103:65:@31.4]
  assign _T_38 = _GEN_0 << 16; // @[Bitwise.scala 103:65:@31.4]
  assign _T_40 = _T_38 & 32'hffff0000; // @[Bitwise.scala 103:75:@33.4]
  assign _T_41 = _T_36 | _T_40; // @[Bitwise.scala 103:39:@34.4]
  assign _T_45 = _T_41[31:8]; // @[Bitwise.scala 103:21:@38.4]
  assign _GEN_1 = {{8'd0}, _T_45}; // @[Bitwise.scala 103:31:@39.4]
  assign _T_46 = _GEN_1 & 32'hff00ff; // @[Bitwise.scala 103:31:@39.4]
  assign _T_47 = _T_41[23:0]; // @[Bitwise.scala 103:46:@40.4]
  assign _GEN_2 = {{8'd0}, _T_47}; // @[Bitwise.scala 103:65:@41.4]
  assign _T_48 = _GEN_2 << 8; // @[Bitwise.scala 103:65:@41.4]
  assign _T_50 = _T_48 & 32'hff00ff00; // @[Bitwise.scala 103:75:@43.4]
  assign _T_51 = _T_46 | _T_50; // @[Bitwise.scala 103:39:@44.4]
  assign _T_55 = _T_51[31:4]; // @[Bitwise.scala 103:21:@48.4]
  assign _GEN_3 = {{4'd0}, _T_55}; // @[Bitwise.scala 103:31:@49.4]
  assign _T_56 = _GEN_3 & 32'hf0f0f0f; // @[Bitwise.scala 103:31:@49.4]
  assign _T_57 = _T_51[27:0]; // @[Bitwise.scala 103:46:@50.4]
  assign _GEN_4 = {{4'd0}, _T_57}; // @[Bitwise.scala 103:65:@51.4]
  assign _T_58 = _GEN_4 << 4; // @[Bitwise.scala 103:65:@51.4]
  assign _T_60 = _T_58 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75:@53.4]
  assign _T_61 = _T_56 | _T_60; // @[Bitwise.scala 103:39:@54.4]
  assign _T_65 = _T_61[31:2]; // @[Bitwise.scala 103:21:@58.4]
  assign _GEN_5 = {{2'd0}, _T_65}; // @[Bitwise.scala 103:31:@59.4]
  assign _T_66 = _GEN_5 & 32'h33333333; // @[Bitwise.scala 103:31:@59.4]
  assign _T_67 = _T_61[29:0]; // @[Bitwise.scala 103:46:@60.4]
  assign _GEN_6 = {{2'd0}, _T_67}; // @[Bitwise.scala 103:65:@61.4]
  assign _T_68 = _GEN_6 << 2; // @[Bitwise.scala 103:65:@61.4]
  assign _T_70 = _T_68 & 32'hcccccccc; // @[Bitwise.scala 103:75:@63.4]
  assign _T_71 = _T_66 | _T_70; // @[Bitwise.scala 103:39:@64.4]
  assign _T_75 = _T_71[31:1]; // @[Bitwise.scala 103:21:@68.4]
  assign _GEN_7 = {{1'd0}, _T_75}; // @[Bitwise.scala 103:31:@69.4]
  assign _T_76 = _GEN_7 & 32'h55555555; // @[Bitwise.scala 103:31:@69.4]
  assign _T_77 = _T_71[30:0]; // @[Bitwise.scala 103:46:@70.4]
  assign _GEN_8 = {{1'd0}, _T_77}; // @[Bitwise.scala 103:65:@71.4]
  assign _T_78 = _GEN_8 << 1; // @[Bitwise.scala 103:65:@71.4]
  assign _T_80 = _T_78 & 32'haaaaaaaa; // @[Bitwise.scala 103:75:@73.4]
  assign _T_81 = _T_76 | _T_80; // @[Bitwise.scala 103:39:@74.4]
  assign shin = _T_30 ? io_A : _T_81; // @[ALU.scala 63:19:@75.4]
  assign _T_83 = shin[31]; // @[ALU.scala 64:41:@77.4]
  assign _T_84 = _T_15 & _T_83; // @[ALU.scala 64:34:@78.4]
  assign _T_85 = {_T_84,shin}; // @[Cat.scala 30:58:@79.4]
  assign _T_86 = $signed(_T_85); // @[ALU.scala 64:57:@80.4]
  assign _T_87 = $signed(_T_86) >>> shamt; // @[ALU.scala 64:64:@81.4]
  assign shiftr = _T_87[31:0]; // @[ALU.scala 64:73:@82.4]
  assign _T_92 = shiftr[31:16]; // @[Bitwise.scala 103:21:@85.4]
  assign _T_93 = {{16'd0}, _T_92}; // @[Bitwise.scala 103:31:@86.4]
  assign _T_94 = shiftr[15:0]; // @[Bitwise.scala 103:46:@87.4]
  assign _GEN_9 = {{16'd0}, _T_94}; // @[Bitwise.scala 103:65:@88.4]
  assign _T_95 = _GEN_9 << 16; // @[Bitwise.scala 103:65:@88.4]
  assign _T_97 = _T_95 & 32'hffff0000; // @[Bitwise.scala 103:75:@90.4]
  assign _T_98 = _T_93 | _T_97; // @[Bitwise.scala 103:39:@91.4]
  assign _T_102 = _T_98[31:8]; // @[Bitwise.scala 103:21:@95.4]
  assign _GEN_10 = {{8'd0}, _T_102}; // @[Bitwise.scala 103:31:@96.4]
  assign _T_103 = _GEN_10 & 32'hff00ff; // @[Bitwise.scala 103:31:@96.4]
  assign _T_104 = _T_98[23:0]; // @[Bitwise.scala 103:46:@97.4]
  assign _GEN_11 = {{8'd0}, _T_104}; // @[Bitwise.scala 103:65:@98.4]
  assign _T_105 = _GEN_11 << 8; // @[Bitwise.scala 103:65:@98.4]
  assign _T_107 = _T_105 & 32'hff00ff00; // @[Bitwise.scala 103:75:@100.4]
  assign _T_108 = _T_103 | _T_107; // @[Bitwise.scala 103:39:@101.4]
  assign _T_112 = _T_108[31:4]; // @[Bitwise.scala 103:21:@105.4]
  assign _GEN_12 = {{4'd0}, _T_112}; // @[Bitwise.scala 103:31:@106.4]
  assign _T_113 = _GEN_12 & 32'hf0f0f0f; // @[Bitwise.scala 103:31:@106.4]
  assign _T_114 = _T_108[27:0]; // @[Bitwise.scala 103:46:@107.4]
  assign _GEN_13 = {{4'd0}, _T_114}; // @[Bitwise.scala 103:65:@108.4]
  assign _T_115 = _GEN_13 << 4; // @[Bitwise.scala 103:65:@108.4]
  assign _T_117 = _T_115 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75:@110.4]
  assign _T_118 = _T_113 | _T_117; // @[Bitwise.scala 103:39:@111.4]
  assign _T_122 = _T_118[31:2]; // @[Bitwise.scala 103:21:@115.4]
  assign _GEN_14 = {{2'd0}, _T_122}; // @[Bitwise.scala 103:31:@116.4]
  assign _T_123 = _GEN_14 & 32'h33333333; // @[Bitwise.scala 103:31:@116.4]
  assign _T_124 = _T_118[29:0]; // @[Bitwise.scala 103:46:@117.4]
  assign _GEN_15 = {{2'd0}, _T_124}; // @[Bitwise.scala 103:65:@118.4]
  assign _T_125 = _GEN_15 << 2; // @[Bitwise.scala 103:65:@118.4]
  assign _T_127 = _T_125 & 32'hcccccccc; // @[Bitwise.scala 103:75:@120.4]
  assign _T_128 = _T_123 | _T_127; // @[Bitwise.scala 103:39:@121.4]
  assign _T_132 = _T_128[31:1]; // @[Bitwise.scala 103:21:@125.4]
  assign _GEN_16 = {{1'd0}, _T_132}; // @[Bitwise.scala 103:31:@126.4]
  assign _T_133 = _GEN_16 & 32'h55555555; // @[Bitwise.scala 103:31:@126.4]
  assign _T_134 = _T_128[30:0]; // @[Bitwise.scala 103:46:@127.4]
  assign _GEN_17 = {{1'd0}, _T_134}; // @[Bitwise.scala 103:65:@128.4]
  assign _T_135 = _GEN_17 << 1; // @[Bitwise.scala 103:65:@128.4]
  assign _T_137 = _T_135 & 32'haaaaaaaa; // @[Bitwise.scala 103:75:@130.4]
  assign shiftl = _T_133 | _T_137; // @[Bitwise.scala 103:39:@131.4]
  assign _T_151 = io_alu_op == 4'h0; // @[ALU.scala 68:19:@132.4]
  assign _T_152 = io_alu_op == 4'h1; // @[ALU.scala 68:44:@133.4]
  assign _T_153 = _T_151 | _T_152; // @[ALU.scala 68:31:@134.4]
  assign _T_154 = io_alu_op == 4'h5; // @[ALU.scala 69:19:@135.4]
  assign _T_155 = io_alu_op == 4'h7; // @[ALU.scala 69:44:@136.4]
  assign _T_156 = _T_154 | _T_155; // @[ALU.scala 69:31:@137.4]
  assign _T_157 = io_alu_op == 4'h9; // @[ALU.scala 70:19:@138.4]
  assign _T_158 = io_alu_op == 4'h8; // @[ALU.scala 70:44:@139.4]
  assign _T_159 = _T_157 | _T_158; // @[ALU.scala 70:31:@140.4]
  assign _T_160 = io_alu_op == 4'h6; // @[ALU.scala 71:19:@141.4]
  assign _T_161 = io_alu_op == 4'h2; // @[ALU.scala 72:19:@142.4]
  assign _T_162 = io_A & io_B; // @[ALU.scala 72:38:@143.4]
  assign _T_163 = io_alu_op == 4'h3; // @[ALU.scala 73:19:@144.4]
  assign _T_164 = io_A | io_B; // @[ALU.scala 73:38:@145.4]
  assign _T_165 = io_alu_op == 4'h4; // @[ALU.scala 74:19:@146.4]
  assign _T_166 = io_A ^ io_B; // @[ALU.scala 74:38:@147.4]
  assign _T_167 = io_alu_op == 4'ha; // @[ALU.scala 75:19:@148.4]
  assign _T_168 = _T_167 ? io_A : io_B; // @[ALU.scala 75:8:@149.4]
  assign _T_169 = _T_165 ? _T_166 : _T_168; // @[ALU.scala 74:8:@150.4]
  assign _T_170 = _T_163 ? _T_164 : _T_169; // @[ALU.scala 73:8:@151.4]
  assign _T_171 = _T_161 ? _T_162 : _T_170; // @[ALU.scala 72:8:@152.4]
  assign _T_172 = _T_160 ? shiftl : _T_171; // @[ALU.scala 71:8:@153.4]
  assign _T_173 = _T_159 ? shiftr : _T_172; // @[ALU.scala 70:8:@154.4]
  assign _T_174 = _T_156 ? {{31'd0}, cmp} : _T_173; // @[ALU.scala 69:8:@155.4]
  assign out = _T_153 ? sum : _T_174; // @[ALU.scala 68:8:@156.4]
  assign io_out = out;
  assign io_sum = sum;
endmodule
module Control( // @[:@160.2]
  input  [31:0] io_inst, // @[:@163.4]
  output [3:0]  io_alu_op // @[:@163.4]
);
  wire [31:0] _T_75; // @[Lookup.scala 9:38:@165.4]
  wire  _T_76; // @[Lookup.scala 9:38:@166.4]
  wire  _T_80; // @[Lookup.scala 9:38:@168.4]
  wire  _T_84; // @[Lookup.scala 9:38:@170.4]
  wire [31:0] _T_87; // @[Lookup.scala 9:38:@171.4]
  wire  _T_88; // @[Lookup.scala 9:38:@172.4]
  wire  _T_92; // @[Lookup.scala 9:38:@174.4]
  wire  _T_96; // @[Lookup.scala 9:38:@176.4]
  wire  _T_100; // @[Lookup.scala 9:38:@178.4]
  wire  _T_104; // @[Lookup.scala 9:38:@180.4]
  wire  _T_108; // @[Lookup.scala 9:38:@182.4]
  wire  _T_112; // @[Lookup.scala 9:38:@184.4]
  wire  _T_116; // @[Lookup.scala 9:38:@186.4]
  wire  _T_120; // @[Lookup.scala 9:38:@188.4]
  wire  _T_124; // @[Lookup.scala 9:38:@190.4]
  wire  _T_128; // @[Lookup.scala 9:38:@192.4]
  wire  _T_132; // @[Lookup.scala 9:38:@194.4]
  wire  _T_136; // @[Lookup.scala 9:38:@196.4]
  wire  _T_140; // @[Lookup.scala 9:38:@198.4]
  wire  _T_144; // @[Lookup.scala 9:38:@200.4]
  wire  _T_148; // @[Lookup.scala 9:38:@202.4]
  wire  _T_152; // @[Lookup.scala 9:38:@204.4]
  wire  _T_156; // @[Lookup.scala 9:38:@206.4]
  wire  _T_160; // @[Lookup.scala 9:38:@208.4]
  wire  _T_164; // @[Lookup.scala 9:38:@210.4]
  wire  _T_168; // @[Lookup.scala 9:38:@212.4]
  wire [31:0] _T_171; // @[Lookup.scala 9:38:@213.4]
  wire  _T_172; // @[Lookup.scala 9:38:@214.4]
  wire  _T_176; // @[Lookup.scala 9:38:@216.4]
  wire  _T_180; // @[Lookup.scala 9:38:@218.4]
  wire  _T_184; // @[Lookup.scala 9:38:@220.4]
  wire  _T_188; // @[Lookup.scala 9:38:@222.4]
  wire  _T_192; // @[Lookup.scala 9:38:@224.4]
  wire  _T_196; // @[Lookup.scala 9:38:@226.4]
  wire  _T_200; // @[Lookup.scala 9:38:@228.4]
  wire  _T_204; // @[Lookup.scala 9:38:@230.4]
  wire  _T_208; // @[Lookup.scala 9:38:@232.4]
  wire  _T_212; // @[Lookup.scala 9:38:@234.4]
  wire  _T_216; // @[Lookup.scala 9:38:@236.4]
  wire  _T_220; // @[Lookup.scala 9:38:@238.4]
  wire [31:0] _T_223; // @[Lookup.scala 9:38:@239.4]
  wire  _T_224; // @[Lookup.scala 9:38:@240.4]
  wire  _T_228; // @[Lookup.scala 9:38:@242.4]
  wire  _T_232; // @[Lookup.scala 9:38:@244.4]
  wire  _T_236; // @[Lookup.scala 9:38:@246.4]
  wire  _T_240; // @[Lookup.scala 9:38:@248.4]
  wire [3:0] _T_468; // @[Lookup.scala 11:37:@466.4]
  wire [3:0] _T_469; // @[Lookup.scala 11:37:@467.4]
  wire [3:0] _T_470; // @[Lookup.scala 11:37:@468.4]
  wire [3:0] _T_471; // @[Lookup.scala 11:37:@469.4]
  wire [3:0] _T_472; // @[Lookup.scala 11:37:@470.4]
  wire [3:0] _T_473; // @[Lookup.scala 11:37:@471.4]
  wire [3:0] _T_474; // @[Lookup.scala 11:37:@472.4]
  wire [3:0] _T_475; // @[Lookup.scala 11:37:@473.4]
  wire [3:0] _T_476; // @[Lookup.scala 11:37:@474.4]
  wire [3:0] _T_477; // @[Lookup.scala 11:37:@475.4]
  wire [3:0] _T_478; // @[Lookup.scala 11:37:@476.4]
  wire [3:0] _T_479; // @[Lookup.scala 11:37:@477.4]
  wire [3:0] _T_480; // @[Lookup.scala 11:37:@478.4]
  wire [3:0] _T_481; // @[Lookup.scala 11:37:@479.4]
  wire [3:0] _T_482; // @[Lookup.scala 11:37:@480.4]
  wire [3:0] _T_483; // @[Lookup.scala 11:37:@481.4]
  wire [3:0] _T_484; // @[Lookup.scala 11:37:@482.4]
  wire [3:0] _T_485; // @[Lookup.scala 11:37:@483.4]
  wire [3:0] _T_486; // @[Lookup.scala 11:37:@484.4]
  wire [3:0] _T_487; // @[Lookup.scala 11:37:@485.4]
  wire [3:0] _T_488; // @[Lookup.scala 11:37:@486.4]
  wire [3:0] _T_489; // @[Lookup.scala 11:37:@487.4]
  wire [3:0] _T_490; // @[Lookup.scala 11:37:@488.4]
  wire [3:0] _T_491; // @[Lookup.scala 11:37:@489.4]
  wire [3:0] _T_492; // @[Lookup.scala 11:37:@490.4]
  wire [3:0] _T_493; // @[Lookup.scala 11:37:@491.4]
  wire [3:0] _T_494; // @[Lookup.scala 11:37:@492.4]
  wire [3:0] _T_495; // @[Lookup.scala 11:37:@493.4]
  wire [3:0] _T_496; // @[Lookup.scala 11:37:@494.4]
  wire [3:0] _T_497; // @[Lookup.scala 11:37:@495.4]
  wire [3:0] _T_498; // @[Lookup.scala 11:37:@496.4]
  wire [3:0] _T_499; // @[Lookup.scala 11:37:@497.4]
  wire [3:0] _T_500; // @[Lookup.scala 11:37:@498.4]
  wire [3:0] _T_501; // @[Lookup.scala 11:37:@499.4]
  wire [3:0] _T_502; // @[Lookup.scala 11:37:@500.4]
  wire [3:0] _T_503; // @[Lookup.scala 11:37:@501.4]
  wire [3:0] _T_504; // @[Lookup.scala 11:37:@502.4]
  wire [3:0] _T_505; // @[Lookup.scala 11:37:@503.4]
  wire [3:0] _T_506; // @[Lookup.scala 11:37:@504.4]
  wire [3:0] _T_507; // @[Lookup.scala 11:37:@505.4]
  wire [3:0] _T_508; // @[Lookup.scala 11:37:@506.4]
  wire [3:0] ctrlSignals_4; // @[Lookup.scala 11:37:@507.4]
  assign _T_75 = io_inst & 32'h7f; // @[Lookup.scala 9:38:@165.4]
  assign _T_76 = 32'h37 == _T_75; // @[Lookup.scala 9:38:@166.4]
  assign _T_80 = 32'h17 == _T_75; // @[Lookup.scala 9:38:@168.4]
  assign _T_84 = 32'h6f == _T_75; // @[Lookup.scala 9:38:@170.4]
  assign _T_87 = io_inst & 32'h707f; // @[Lookup.scala 9:38:@171.4]
  assign _T_88 = 32'h67 == _T_87; // @[Lookup.scala 9:38:@172.4]
  assign _T_92 = 32'h63 == _T_87; // @[Lookup.scala 9:38:@174.4]
  assign _T_96 = 32'h1063 == _T_87; // @[Lookup.scala 9:38:@176.4]
  assign _T_100 = 32'h4063 == _T_87; // @[Lookup.scala 9:38:@178.4]
  assign _T_104 = 32'h5063 == _T_87; // @[Lookup.scala 9:38:@180.4]
  assign _T_108 = 32'h6063 == _T_87; // @[Lookup.scala 9:38:@182.4]
  assign _T_112 = 32'h7063 == _T_87; // @[Lookup.scala 9:38:@184.4]
  assign _T_116 = 32'h3 == _T_87; // @[Lookup.scala 9:38:@186.4]
  assign _T_120 = 32'h1003 == _T_87; // @[Lookup.scala 9:38:@188.4]
  assign _T_124 = 32'h2003 == _T_87; // @[Lookup.scala 9:38:@190.4]
  assign _T_128 = 32'h4003 == _T_87; // @[Lookup.scala 9:38:@192.4]
  assign _T_132 = 32'h5003 == _T_87; // @[Lookup.scala 9:38:@194.4]
  assign _T_136 = 32'h23 == _T_87; // @[Lookup.scala 9:38:@196.4]
  assign _T_140 = 32'h1023 == _T_87; // @[Lookup.scala 9:38:@198.4]
  assign _T_144 = 32'h2023 == _T_87; // @[Lookup.scala 9:38:@200.4]
  assign _T_148 = 32'h13 == _T_87; // @[Lookup.scala 9:38:@202.4]
  assign _T_152 = 32'h2013 == _T_87; // @[Lookup.scala 9:38:@204.4]
  assign _T_156 = 32'h3013 == _T_87; // @[Lookup.scala 9:38:@206.4]
  assign _T_160 = 32'h4013 == _T_87; // @[Lookup.scala 9:38:@208.4]
  assign _T_164 = 32'h6013 == _T_87; // @[Lookup.scala 9:38:@210.4]
  assign _T_168 = 32'h7013 == _T_87; // @[Lookup.scala 9:38:@212.4]
  assign _T_171 = io_inst & 32'hfe00707f; // @[Lookup.scala 9:38:@213.4]
  assign _T_172 = 32'h1013 == _T_171; // @[Lookup.scala 9:38:@214.4]
  assign _T_176 = 32'h5013 == _T_171; // @[Lookup.scala 9:38:@216.4]
  assign _T_180 = 32'h40005013 == _T_171; // @[Lookup.scala 9:38:@218.4]
  assign _T_184 = 32'h33 == _T_171; // @[Lookup.scala 9:38:@220.4]
  assign _T_188 = 32'h40000033 == _T_171; // @[Lookup.scala 9:38:@222.4]
  assign _T_192 = 32'h1033 == _T_171; // @[Lookup.scala 9:38:@224.4]
  assign _T_196 = 32'h2033 == _T_171; // @[Lookup.scala 9:38:@226.4]
  assign _T_200 = 32'h3033 == _T_171; // @[Lookup.scala 9:38:@228.4]
  assign _T_204 = 32'h4033 == _T_171; // @[Lookup.scala 9:38:@230.4]
  assign _T_208 = 32'h5033 == _T_171; // @[Lookup.scala 9:38:@232.4]
  assign _T_212 = 32'h40005033 == _T_171; // @[Lookup.scala 9:38:@234.4]
  assign _T_216 = 32'h6033 == _T_171; // @[Lookup.scala 9:38:@236.4]
  assign _T_220 = 32'h7033 == _T_171; // @[Lookup.scala 9:38:@238.4]
  assign _T_223 = io_inst & 32'hf00fffff; // @[Lookup.scala 9:38:@239.4]
  assign _T_224 = 32'hf == _T_223; // @[Lookup.scala 9:38:@240.4]
  assign _T_228 = 32'h100f == io_inst; // @[Lookup.scala 9:38:@242.4]
  assign _T_232 = 32'h1073 == _T_87; // @[Lookup.scala 9:38:@244.4]
  assign _T_236 = 32'h2073 == _T_87; // @[Lookup.scala 9:38:@246.4]
  assign _T_240 = 32'h3073 == _T_87; // @[Lookup.scala 9:38:@248.4]
  assign _T_468 = _T_240 ? 4'ha : 4'hf; // @[Lookup.scala 11:37:@466.4]
  assign _T_469 = _T_236 ? 4'ha : _T_468; // @[Lookup.scala 11:37:@467.4]
  assign _T_470 = _T_232 ? 4'ha : _T_469; // @[Lookup.scala 11:37:@468.4]
  assign _T_471 = _T_228 ? 4'hf : _T_470; // @[Lookup.scala 11:37:@469.4]
  assign _T_472 = _T_224 ? 4'hf : _T_471; // @[Lookup.scala 11:37:@470.4]
  assign _T_473 = _T_220 ? 4'h2 : _T_472; // @[Lookup.scala 11:37:@471.4]
  assign _T_474 = _T_216 ? 4'h3 : _T_473; // @[Lookup.scala 11:37:@472.4]
  assign _T_475 = _T_212 ? 4'h9 : _T_474; // @[Lookup.scala 11:37:@473.4]
  assign _T_476 = _T_208 ? 4'h8 : _T_475; // @[Lookup.scala 11:37:@474.4]
  assign _T_477 = _T_204 ? 4'h4 : _T_476; // @[Lookup.scala 11:37:@475.4]
  assign _T_478 = _T_200 ? 4'h7 : _T_477; // @[Lookup.scala 11:37:@476.4]
  assign _T_479 = _T_196 ? 4'h5 : _T_478; // @[Lookup.scala 11:37:@477.4]
  assign _T_480 = _T_192 ? 4'h6 : _T_479; // @[Lookup.scala 11:37:@478.4]
  assign _T_481 = _T_188 ? 4'h1 : _T_480; // @[Lookup.scala 11:37:@479.4]
  assign _T_482 = _T_184 ? 4'h0 : _T_481; // @[Lookup.scala 11:37:@480.4]
  assign _T_483 = _T_180 ? 4'h9 : _T_482; // @[Lookup.scala 11:37:@481.4]
  assign _T_484 = _T_176 ? 4'h8 : _T_483; // @[Lookup.scala 11:37:@482.4]
  assign _T_485 = _T_172 ? 4'h6 : _T_484; // @[Lookup.scala 11:37:@483.4]
  assign _T_486 = _T_168 ? 4'h2 : _T_485; // @[Lookup.scala 11:37:@484.4]
  assign _T_487 = _T_164 ? 4'h3 : _T_486; // @[Lookup.scala 11:37:@485.4]
  assign _T_488 = _T_160 ? 4'h4 : _T_487; // @[Lookup.scala 11:37:@486.4]
  assign _T_489 = _T_156 ? 4'h7 : _T_488; // @[Lookup.scala 11:37:@487.4]
  assign _T_490 = _T_152 ? 4'h5 : _T_489; // @[Lookup.scala 11:37:@488.4]
  assign _T_491 = _T_148 ? 4'h0 : _T_490; // @[Lookup.scala 11:37:@489.4]
  assign _T_492 = _T_144 ? 4'h0 : _T_491; // @[Lookup.scala 11:37:@490.4]
  assign _T_493 = _T_140 ? 4'h0 : _T_492; // @[Lookup.scala 11:37:@491.4]
  assign _T_494 = _T_136 ? 4'h0 : _T_493; // @[Lookup.scala 11:37:@492.4]
  assign _T_495 = _T_132 ? 4'h0 : _T_494; // @[Lookup.scala 11:37:@493.4]
  assign _T_496 = _T_128 ? 4'h0 : _T_495; // @[Lookup.scala 11:37:@494.4]
  assign _T_497 = _T_124 ? 4'h0 : _T_496; // @[Lookup.scala 11:37:@495.4]
  assign _T_498 = _T_120 ? 4'h0 : _T_497; // @[Lookup.scala 11:37:@496.4]
  assign _T_499 = _T_116 ? 4'h0 : _T_498; // @[Lookup.scala 11:37:@497.4]
  assign _T_500 = _T_112 ? 4'h0 : _T_499; // @[Lookup.scala 11:37:@498.4]
  assign _T_501 = _T_108 ? 4'h0 : _T_500; // @[Lookup.scala 11:37:@499.4]
  assign _T_502 = _T_104 ? 4'h0 : _T_501; // @[Lookup.scala 11:37:@500.4]
  assign _T_503 = _T_100 ? 4'h0 : _T_502; // @[Lookup.scala 11:37:@501.4]
  assign _T_504 = _T_96 ? 4'h0 : _T_503; // @[Lookup.scala 11:37:@502.4]
  assign _T_505 = _T_92 ? 4'h0 : _T_504; // @[Lookup.scala 11:37:@503.4]
  assign _T_506 = _T_88 ? 4'h0 : _T_505; // @[Lookup.scala 11:37:@504.4]
  assign _T_507 = _T_84 ? 4'h0 : _T_506; // @[Lookup.scala 11:37:@505.4]
  assign _T_508 = _T_80 ? 4'h0 : _T_507; // @[Lookup.scala 11:37:@506.4]
  assign ctrlSignals_4 = _T_76 ? 4'hb : _T_508; // @[Lookup.scala 11:37:@507.4]
  assign io_alu_op = ctrlSignals_4;
endmodule
module ALUTester( // @[:@916.2]
  input   clock, // @[:@917.4]
  input   reset // @[:@918.4]
);
  wire [31:0] dut_io_A; // @[ALUTests.scala 11:19:@921.4]
  wire [31:0] dut_io_B; // @[ALUTests.scala 11:19:@921.4]
  wire [3:0] dut_io_alu_op; // @[ALUTests.scala 11:19:@921.4]
  wire [31:0] dut_io_out; // @[ALUTests.scala 11:19:@921.4]
  wire [31:0] dut_io_sum; // @[ALUTests.scala 11:19:@921.4]
  wire [31:0] ctrl_io_inst; // @[ALUTests.scala 12:20:@924.4]
  wire [3:0] ctrl_io_alu_op; // @[ALUTests.scala 12:20:@924.4]
  reg [5:0] value; // @[Counter.scala 26:33:@927.4]
  reg [31:0] _RAND_0;
  wire  done; // @[Counter.scala 34:24:@929.6]
  wire [6:0] _T_610; // @[Counter.scala 35:22:@930.6]
  wire [5:0] _T_611; // @[Counter.scala 35:22:@931.6]
  wire [5:0] _GEN_0; // @[Counter.scala 37:21:@933.6]
  wire  _T_1653; // @[ALUTests.scala 28:32:@1448.4]
  wire  _T_1655; // @[ALUTests.scala 29:32:@1449.4]
  wire  _T_1657; // @[ALUTests.scala 30:32:@1450.4]
  wire  _T_1659; // @[ALUTests.scala 31:32:@1451.4]
  wire  _T_1661; // @[ALUTests.scala 32:32:@1452.4]
  wire  _T_1663; // @[ALUTests.scala 33:32:@1453.4]
  wire  _T_1665; // @[ALUTests.scala 34:32:@1454.4]
  wire  _T_1667; // @[ALUTests.scala 35:32:@1455.4]
  wire  _T_1669; // @[ALUTests.scala 36:32:@1456.4]
  wire  _T_1671; // @[ALUTests.scala 37:32:@1457.4]
  wire  _T_1673; // @[ALUTests.scala 38:32:@1458.4]
  wire [31:0] _T_1674; // @[ALUTests.scala 38:17:@1459.4]
  wire [31:0] _GEN_3; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_4; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_5; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_6; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_7; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_8; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_9; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_10; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_11; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_12; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_13; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_14; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_15; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_16; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_17; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_18; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_19; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_20; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_21; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_22; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_23; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_24; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_25; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_26; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_27; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_28; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_29; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_30; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_31; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_32; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_33; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_34; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_35; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_36; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_37; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_38; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_39; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_40; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_41; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_42; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_43; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_44; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_45; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_46; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_47; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_48; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_49; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_50; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_51; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _T_1675; // @[ALUTests.scala 37:17:@1460.4]
  wire [31:0] _GEN_53; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_54; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_55; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_56; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_57; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_58; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_59; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_60; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_61; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_62; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_63; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_64; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_65; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_66; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_67; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_68; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_69; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_70; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_71; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_72; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_73; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_74; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_75; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_76; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_77; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_78; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_79; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_80; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_81; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_82; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_83; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_84; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_85; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_86; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_87; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_88; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_89; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_90; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_91; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_92; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_93; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_94; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_95; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_96; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_97; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_98; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_99; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_100; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_101; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _T_1676; // @[ALUTests.scala 36:17:@1461.4]
  wire [31:0] _GEN_103; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_104; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_105; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_106; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_107; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_108; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_109; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_110; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_111; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_112; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_113; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_114; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_115; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_116; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_117; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_118; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_119; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_120; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_121; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_122; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_123; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_124; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_125; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_126; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_127; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_128; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_129; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_130; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_131; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_132; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_133; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_134; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_135; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_136; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_137; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_138; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_139; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_140; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_141; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_142; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_143; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_144; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_145; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_146; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_147; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_148; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_149; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_150; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_151; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _T_1677; // @[ALUTests.scala 35:17:@1462.4]
  wire [31:0] _GEN_154; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_155; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_156; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_157; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_158; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_159; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_160; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_161; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_162; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_163; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_164; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_165; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_166; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_167; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_168; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_169; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_170; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_171; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_172; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_173; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_174; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_175; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_176; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_177; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_178; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_179; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_180; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_181; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_182; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_183; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_184; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_185; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_186; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_187; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_188; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_189; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_190; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_191; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_192; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_193; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_194; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_195; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_196; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_197; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_198; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_199; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_200; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_201; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _T_1678; // @[ALUTests.scala 34:17:@1463.4]
  wire [31:0] _GEN_203; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_204; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_205; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_206; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_207; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_208; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_209; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_210; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_211; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_212; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_213; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_214; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_215; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_216; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_217; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_218; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_219; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_220; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_221; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_222; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_223; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_224; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_225; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_226; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_227; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_228; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_229; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_230; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_231; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_232; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_233; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_234; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_235; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_236; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_237; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_238; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_239; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_240; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_241; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_242; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_243; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_244; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_245; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_246; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_247; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_248; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_249; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_250; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_251; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _T_1679; // @[ALUTests.scala 33:17:@1464.4]
  wire [31:0] _GEN_253; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_254; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_255; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_256; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_257; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_258; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_259; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_260; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_261; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_262; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_263; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_264; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_265; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_266; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_267; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_268; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_269; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_270; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_271; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_272; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_273; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_274; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_275; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_276; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_277; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_278; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_279; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_280; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_281; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_282; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_283; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_284; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_285; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_286; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_287; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_288; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_289; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_290; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_291; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_292; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_293; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_294; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_295; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_296; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_297; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_298; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_299; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_300; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_301; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _T_1680; // @[ALUTests.scala 32:17:@1465.4]
  wire [31:0] _GEN_303; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_304; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_305; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_306; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_307; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_308; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_309; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_310; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_311; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_312; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_313; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_314; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_315; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_316; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_317; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_318; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_319; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_320; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_321; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_322; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_323; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_324; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_325; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_326; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_327; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_328; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_329; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_330; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_331; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_332; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_333; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_334; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_335; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_336; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_337; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_338; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_339; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_340; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_341; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_342; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_343; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_344; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_345; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_346; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_347; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_348; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_349; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_350; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_351; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _T_1681; // @[ALUTests.scala 31:17:@1466.4]
  wire [31:0] _GEN_353; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_354; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_355; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_356; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_357; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_358; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_359; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_360; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_361; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_362; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_363; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_364; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_365; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_366; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_367; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_368; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_369; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_370; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_371; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_372; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_373; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_374; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_375; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_376; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_377; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_378; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_379; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_380; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_381; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_382; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_383; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_384; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_385; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_386; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_387; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_388; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_389; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_390; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_391; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_392; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_393; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_394; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_395; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_396; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_397; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_398; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_399; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_400; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_401; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _T_1682; // @[ALUTests.scala 30:17:@1467.4]
  wire [31:0] _GEN_403; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_404; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_405; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_406; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_407; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_408; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_409; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_410; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_411; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_412; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_413; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_414; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_415; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_416; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_417; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_418; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_419; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_420; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_421; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_422; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_423; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_424; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_425; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_426; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_427; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_428; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_429; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_430; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_431; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_432; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_433; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_434; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_435; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_436; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_437; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_438; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_439; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_440; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_441; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_442; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_443; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_444; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_445; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_446; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_447; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_448; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_449; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_450; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_451; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _T_1683; // @[ALUTests.scala 29:17:@1468.4]
  wire [31:0] _GEN_453; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_454; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_455; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_456; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_457; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_458; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_459; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_460; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_461; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_462; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_463; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_464; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_465; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_466; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_467; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_468; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_469; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_470; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_471; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_472; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_473; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_474; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_475; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_476; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_477; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_478; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_479; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_480; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_481; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_482; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_483; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_484; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_485; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_486; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_487; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_488; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_489; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_490; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_491; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_492; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_493; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_494; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_495; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_496; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_497; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_498; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_499; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_500; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _GEN_501; // @[ALUTests.scala 28:17:@1469.4]
  wire [31:0] _T_1684; // @[ALUTests.scala 28:17:@1469.4]
  wire  _T_1685; // @[ALUTests.scala 39:31:@1470.4]
  wire [31:0] _T_1688; // @[ALUTests.scala 39:17:@1471.4]
  wire [31:0] _GEN_503; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_504; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_505; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_506; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_507; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_508; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_509; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_510; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_511; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_512; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_513; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_514; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_515; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_516; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_517; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_518; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_519; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_520; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_521; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_522; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_523; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_524; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_525; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_526; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_527; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_528; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_529; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_530; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_531; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_532; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_533; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_534; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_535; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_536; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_537; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_538; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_539; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_540; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_541; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_542; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_543; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_544; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_545; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_546; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_547; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_548; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_549; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_550; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_551; // @[ALUTests.scala 41:16:@1523.4]
  wire [31:0] _GEN_553; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_554; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_555; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_556; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_557; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_558; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_559; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_560; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_561; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_562; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_563; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_564; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_565; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_566; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_567; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_568; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_569; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_570; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_571; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_572; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_573; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_574; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_575; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_576; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_577; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_578; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_579; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_580; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_581; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_582; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_583; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_584; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_585; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_586; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_587; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_588; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_589; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_590; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_591; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_592; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_593; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_594; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_595; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_596; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_597; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_598; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_599; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_600; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_601; // @[ALUTests.scala 43:12:@1576.4]
  wire [31:0] _GEN_603; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_604; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_605; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_606; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_607; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_608; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_609; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_610; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_611; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_612; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_613; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_614; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_615; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_616; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_617; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_618; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_619; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_620; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_621; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_622; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_623; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_624; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_625; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_626; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_627; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_628; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_629; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_630; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_631; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_632; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_633; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_634; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_635; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_636; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_637; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_638; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_639; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_640; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_641; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_642; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_643; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_644; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_645; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_646; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_647; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_648; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_649; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_650; // @[ALUTests.scala 44:12:@1628.4]
  wire [31:0] _GEN_651; // @[ALUTests.scala 44:12:@1628.4]
  wire  _T_1959; // @[ALUTests.scala 46:20:@1631.6]
  wire  _T_1963; // @[ALUTests.scala 47:21:@1641.4]
  wire  _T_1965; // @[ALUTests.scala 47:9:@1643.4]
  wire  _T_1967; // @[ALUTests.scala 47:9:@1644.4]
  wire  _T_1968; // @[ALUTests.scala 48:21:@1649.4]
  wire  _T_1970; // @[ALUTests.scala 48:9:@1651.4]
  wire  _T_1972; // @[ALUTests.scala 48:9:@1652.4]
  ALUArea dut ( // @[ALUTests.scala 11:19:@921.4]
    .io_A(dut_io_A),
    .io_B(dut_io_B),
    .io_alu_op(dut_io_alu_op),
    .io_out(dut_io_out),
    .io_sum(dut_io_sum)
  );
  Control ctrl ( // @[ALUTests.scala 12:20:@924.4]
    .io_inst(ctrl_io_inst),
    .io_alu_op(ctrl_io_alu_op)
  );
  assign done = value == 6'h31; // @[Counter.scala 34:24:@929.6]
  assign _T_610 = value + 6'h1; // @[Counter.scala 35:22:@930.6]
  assign _T_611 = _T_610[5:0]; // @[Counter.scala 35:22:@931.6]
  assign _GEN_0 = done ? 6'h0 : _T_611; // @[Counter.scala 37:21:@933.6]
  assign _T_1653 = dut_io_alu_op == 4'h0; // @[ALUTests.scala 28:32:@1448.4]
  assign _T_1655 = dut_io_alu_op == 4'h1; // @[ALUTests.scala 29:32:@1449.4]
  assign _T_1657 = dut_io_alu_op == 4'h2; // @[ALUTests.scala 30:32:@1450.4]
  assign _T_1659 = dut_io_alu_op == 4'h3; // @[ALUTests.scala 31:32:@1451.4]
  assign _T_1661 = dut_io_alu_op == 4'h4; // @[ALUTests.scala 32:32:@1452.4]
  assign _T_1663 = dut_io_alu_op == 4'h5; // @[ALUTests.scala 33:32:@1453.4]
  assign _T_1665 = dut_io_alu_op == 4'h7; // @[ALUTests.scala 34:32:@1454.4]
  assign _T_1667 = dut_io_alu_op == 4'h6; // @[ALUTests.scala 35:32:@1455.4]
  assign _T_1669 = dut_io_alu_op == 4'h8; // @[ALUTests.scala 36:32:@1456.4]
  assign _T_1671 = dut_io_alu_op == 4'h9; // @[ALUTests.scala 37:32:@1457.4]
  assign _T_1673 = dut_io_alu_op == 4'ha; // @[ALUTests.scala 38:32:@1458.4]
  assign _T_1674 = _T_1673 ? dut_io_A : dut_io_B; // @[ALUTests.scala 38:17:@1459.4]
  assign _GEN_3 = 6'h1 == value ? 32'h3f8888c : 32'hffffffca; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_4 = 6'h2 == value ? 32'hffffffd5 : _GEN_3; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_5 = 6'h3 == value ? 32'h3b4a9 : _GEN_4; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_6 = 6'h4 == value ? 32'h3c6bbbf : _GEN_5; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_7 = 6'h5 == value ? 32'h69c : _GEN_6; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_8 = 6'h6 == value ? 32'h90 : _GEN_7; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_9 = 6'h7 == value ? 32'hb03 : _GEN_8; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_10 = 6'h8 == value ? 32'hffffff43 : _GEN_9; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_11 = 6'h9 == value ? 32'h1199b : _GEN_10; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_12 = 6'ha == value ? 32'hffcd8fa0 : _GEN_11; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_13 = 6'hb == value ? 32'hffffc4bc : _GEN_12; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_14 = 6'hc == value ? 32'h143 : _GEN_13; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_15 = 6'hd == value ? 32'h1da58d03 : _GEN_14; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_16 = 6'he == value ? 32'hbab34d5 : _GEN_15; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_17 = 6'hf == value ? 32'h15 : _GEN_16; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_18 = 6'h10 == value ? 32'h74 : _GEN_17; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_19 = 6'h11 == value ? 32'hffffffed : _GEN_18; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_20 = 6'h12 == value ? 32'h11054e26 : _GEN_19; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_21 = 6'h13 == value ? 32'hfffffff9 : _GEN_20; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_22 = 6'h14 == value ? 32'h4 : _GEN_21; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_23 = 6'h15 == value ? 32'hffffffa0 : _GEN_22; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_24 = 6'h16 == value ? 32'h0 : _GEN_23; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_25 = 6'h17 == value ? 32'hffffffaf : _GEN_24; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_26 = 6'h18 == value ? 32'hfffffffb : _GEN_25; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_27 = 6'h19 == value ? 32'h774a : _GEN_26; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_28 = 6'h1a == value ? 32'h3eb71fbf : _GEN_27; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_29 = 6'h1b == value ? 32'hffffffb2 : _GEN_28; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_30 = 6'h1c == value ? 32'h1d51 : _GEN_29; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_31 = 6'h1d == value ? 32'hfffff93d : _GEN_30; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_32 = 6'h1e == value ? 32'hfffff3bc : _GEN_31; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_33 = 6'h1f == value ? 32'hffffffff : _GEN_32; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_34 = 6'h20 == value ? 32'he4827569 : _GEN_33; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_35 = 6'h21 == value ? 32'hfd76a50b : _GEN_34; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_36 = 6'h22 == value ? 32'hffffff9d : _GEN_35; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_37 = 6'h23 == value ? 32'h2 : _GEN_36; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_38 = 6'h24 == value ? 32'he7986f : _GEN_37; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_39 = 6'h25 == value ? 32'h358 : _GEN_38; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_40 = 6'h26 == value ? 32'hffffffd6 : _GEN_39; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_41 = 6'h27 == value ? 32'h10fcdd0 : _GEN_40; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_42 = 6'h28 == value ? 32'hffffd2c7 : _GEN_41; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_43 = 6'h29 == value ? 32'hffc63482 : _GEN_42; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_44 = 6'h2a == value ? 32'hffd13a9f : _GEN_43; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_45 = 6'h2b == value ? 32'he87d8226 : _GEN_44; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_46 = 6'h2c == value ? 32'h11983c8 : _GEN_45; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_47 = 6'h2d == value ? 32'h16096fdd : _GEN_46; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_48 = 6'h2e == value ? 32'ha69bb37b : _GEN_47; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_49 = 6'h2f == value ? 32'hff9c12ad : _GEN_48; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_50 = 6'h30 == value ? 32'hfff55c9f : _GEN_49; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_51 = 6'h31 == value ? 32'h6a7 : _GEN_50; // @[ALUTests.scala 37:17:@1460.4]
  assign _T_1675 = _T_1671 ? _GEN_51 : _T_1674; // @[ALUTests.scala 37:17:@1460.4]
  assign _GEN_53 = 6'h1 == value ? 32'h3f8888c : 32'h4a; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_54 = 6'h2 == value ? 32'h55 : _GEN_53; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_55 = 6'h3 == value ? 32'h3b4a9 : _GEN_54; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_56 = 6'h4 == value ? 32'h3c6bbbf : _GEN_55; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_57 = 6'h5 == value ? 32'h69c : _GEN_56; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_58 = 6'h6 == value ? 32'h90 : _GEN_57; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_59 = 6'h7 == value ? 32'hb03 : _GEN_58; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_60 = 6'h8 == value ? 32'h743 : _GEN_59; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_61 = 6'h9 == value ? 32'h1199b : _GEN_60; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_62 = 6'ha == value ? 32'h4d8fa0 : _GEN_61; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_63 = 6'hb == value ? 32'h44bc : _GEN_62; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_64 = 6'hc == value ? 32'h143 : _GEN_63; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_65 = 6'hd == value ? 32'h1da58d03 : _GEN_64; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_66 = 6'he == value ? 32'hbab34d5 : _GEN_65; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_67 = 6'hf == value ? 32'h15 : _GEN_66; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_68 = 6'h10 == value ? 32'h74 : _GEN_67; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_69 = 6'h11 == value ? 32'hed : _GEN_68; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_70 = 6'h12 == value ? 32'h11054e26 : _GEN_69; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_71 = 6'h13 == value ? 32'h39 : _GEN_70; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_72 = 6'h14 == value ? 32'h4 : _GEN_71; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_73 = 6'h15 == value ? 32'ha0 : _GEN_72; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_74 = 6'h16 == value ? 32'h0 : _GEN_73; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_75 = 6'h17 == value ? 32'haf : _GEN_74; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_76 = 6'h18 == value ? 32'hb : _GEN_75; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_77 = 6'h19 == value ? 32'h774a : _GEN_76; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_78 = 6'h1a == value ? 32'h3eb71fbf : _GEN_77; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_79 = 6'h1b == value ? 32'h1b2 : _GEN_78; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_80 = 6'h1c == value ? 32'h1d51 : _GEN_79; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_81 = 6'h1d == value ? 32'h93d : _GEN_80; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_82 = 6'h1e == value ? 32'h13bc : _GEN_81; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_83 = 6'h1f == value ? 32'h1 : _GEN_82; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_84 = 6'h20 == value ? 32'h24827569 : _GEN_83; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_85 = 6'h21 == value ? 32'h576a50b : _GEN_84; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_86 = 6'h22 == value ? 32'h39d : _GEN_85; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_87 = 6'h23 == value ? 32'h2 : _GEN_86; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_88 = 6'h24 == value ? 32'he7986f : _GEN_87; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_89 = 6'h25 == value ? 32'h358 : _GEN_88; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_90 = 6'h26 == value ? 32'h56 : _GEN_89; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_91 = 6'h27 == value ? 32'h10fcdd0 : _GEN_90; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_92 = 6'h28 == value ? 32'h52c7 : _GEN_91; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_93 = 6'h29 == value ? 32'h463482 : _GEN_92; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_94 = 6'h2a == value ? 32'h1d13a9f : _GEN_93; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_95 = 6'h2b == value ? 32'h287d8226 : _GEN_94; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_96 = 6'h2c == value ? 32'h11983c8 : _GEN_95; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_97 = 6'h2d == value ? 32'h16096fdd : _GEN_96; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_98 = 6'h2e == value ? 32'ha69bb37b : _GEN_97; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_99 = 6'h2f == value ? 32'h19c12ad : _GEN_98; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_100 = 6'h30 == value ? 32'h155c9f : _GEN_99; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_101 = 6'h31 == value ? 32'h6a7 : _GEN_100; // @[ALUTests.scala 36:17:@1461.4]
  assign _T_1676 = _T_1669 ? _GEN_101 : _T_1675; // @[ALUTests.scala 36:17:@1461.4]
  assign _GEN_103 = 6'h1 == value ? 32'he2223100 : 32'h4a000000; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_104 = 6'h2 == value ? 32'h3c000000 : _GEN_103; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_105 = 6'h3 == value ? 32'h2a438000 : _GEN_104; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_106 = 6'h4 == value ? 32'hc6bbbf30 : _GEN_105; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_107 = 6'h5 == value ? 32'h8500000 : _GEN_106; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_108 = 6'h6 == value ? 32'h7d000000 : _GEN_107; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_109 = 6'h7 == value ? 32'h33680000 : _GEN_108; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_110 = 6'h8 == value ? 32'h44200000 : _GEN_109; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_111 = 6'h9 == value ? 32'hbd1d8000 : _GEN_110; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_112 = 6'ha == value ? 32'h3e832600 : _GEN_111; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_113 = 6'hb == value ? 32'ha5660000 : _GEN_112; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_114 = 6'hc == value ? 32'hc1000000 : _GEN_113; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_115 = 6'hd == value ? 32'hda58d030 : _GEN_114; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_116 = 6'he == value ? 32'heacd3558 : _GEN_115; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_117 = 6'hf == value ? 32'h4c000000 : _GEN_116; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_118 = 6'h10 == value ? 32'h96200000 : _GEN_117; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_119 = 6'h11 == value ? 32'h2d000000 : _GEN_118; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_120 = 6'h12 == value ? 32'h1054e268 : _GEN_119; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_121 = 6'h13 == value ? 32'ha8000000 : _GEN_120; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_122 = 6'h14 == value ? 32'hb0000000 : _GEN_121; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_123 = 6'h15 == value ? 32'h44000000 : _GEN_122; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_124 = 6'h16 == value ? 32'h80000000 : _GEN_123; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_125 = 6'h17 == value ? 32'ha6000000 : _GEN_124; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_126 = 6'h18 == value ? 32'he0000000 : _GEN_125; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_127 = 6'h19 == value ? 32'h50e30000 : _GEN_126; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_128 = 6'h1a == value ? 32'hfadc7efc : _GEN_127; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_129 = 6'h1b == value ? 32'hc4000000 : _GEN_128; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_130 = 6'h1c == value ? 32'hf50f0000 : _GEN_129; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_131 = 6'h1d == value ? 32'h22c00000 : _GEN_130; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_132 = 6'h1e == value ? 32'h4c080000 : _GEN_131; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_133 = 6'h1f == value ? 32'h80000000 : _GEN_132; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_134 = 6'h20 == value ? 32'h4827569c : _GEN_133; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_135 = 6'h21 == value ? 32'hda942e40 : _GEN_134; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_136 = 6'h22 == value ? 32'h37800000 : _GEN_135; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_137 = 6'h23 == value ? 32'h40000000 : _GEN_136; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_138 = 6'h24 == value ? 32'he61bc380 : _GEN_137; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_139 = 6'h25 == value ? 32'hd1f00000 : _GEN_138; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_140 = 6'h26 == value ? 32'ha000000 : _GEN_139; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_141 = 6'h27 == value ? 32'hfcdd0a80 : _GEN_140; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_142 = 6'h28 == value ? 32'hec3c0000 : _GEN_141; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_143 = 6'h29 == value ? 32'hd20bae00 : _GEN_142; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_144 = 6'h2a == value ? 32'h4ea7d800 : _GEN_143; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_145 = 6'h2b == value ? 32'h87d82264 : _GEN_144; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_146 = 6'h2c == value ? 32'h660f2140 : _GEN_145; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_147 = 6'h2d == value ? 32'h16096fdd : _GEN_146; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_148 = 6'h2e == value ? 32'ha69bb37b : _GEN_147; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_149 = 6'h2f == value ? 32'h4ab5900 : _GEN_148; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_150 = 6'h30 == value ? 32'h27fe5800 : _GEN_149; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_151 = 6'h31 == value ? 32'h6b600000 : _GEN_150; // @[ALUTests.scala 35:17:@1462.4]
  assign _T_1677 = _T_1667 ? _GEN_151 : _T_1676; // @[ALUTests.scala 35:17:@1462.4]
  assign _GEN_154 = 6'h2 == value ? 32'h0 : 32'h1; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_155 = 6'h3 == value ? 32'h1 : _GEN_154; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_156 = 6'h4 == value ? 32'h1 : _GEN_155; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_157 = 6'h5 == value ? 32'h1 : _GEN_156; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_158 = 6'h6 == value ? 32'h1 : _GEN_157; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_159 = 6'h7 == value ? 32'h1 : _GEN_158; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_160 = 6'h8 == value ? 32'h1 : _GEN_159; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_161 = 6'h9 == value ? 32'h1 : _GEN_160; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_162 = 6'ha == value ? 32'h0 : _GEN_161; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_163 = 6'hb == value ? 32'h0 : _GEN_162; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_164 = 6'hc == value ? 32'h1 : _GEN_163; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_165 = 6'hd == value ? 32'h1 : _GEN_164; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_166 = 6'he == value ? 32'h0 : _GEN_165; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_167 = 6'hf == value ? 32'h1 : _GEN_166; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_168 = 6'h10 == value ? 32'h0 : _GEN_167; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_169 = 6'h11 == value ? 32'h0 : _GEN_168; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_170 = 6'h12 == value ? 32'h1 : _GEN_169; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_171 = 6'h13 == value ? 32'h1 : _GEN_170; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_172 = 6'h14 == value ? 32'h1 : _GEN_171; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_173 = 6'h15 == value ? 32'h0 : _GEN_172; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_174 = 6'h16 == value ? 32'h1 : _GEN_173; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_175 = 6'h17 == value ? 32'h1 : _GEN_174; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_176 = 6'h18 == value ? 32'h1 : _GEN_175; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_177 = 6'h19 == value ? 32'h1 : _GEN_176; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_178 = 6'h1a == value ? 32'h0 : _GEN_177; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_179 = 6'h1b == value ? 32'h1 : _GEN_178; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_180 = 6'h1c == value ? 32'h1 : _GEN_179; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_181 = 6'h1d == value ? 32'h0 : _GEN_180; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_182 = 6'h1e == value ? 32'h0 : _GEN_181; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_183 = 6'h1f == value ? 32'h0 : _GEN_182; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_184 = 6'h20 == value ? 32'h1 : _GEN_183; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_185 = 6'h21 == value ? 32'h1 : _GEN_184; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_186 = 6'h22 == value ? 32'h0 : _GEN_185; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_187 = 6'h23 == value ? 32'h1 : _GEN_186; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_188 = 6'h24 == value ? 32'h1 : _GEN_187; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_189 = 6'h25 == value ? 32'h1 : _GEN_188; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_190 = 6'h26 == value ? 32'h1 : _GEN_189; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_191 = 6'h27 == value ? 32'h1 : _GEN_190; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_192 = 6'h28 == value ? 32'h0 : _GEN_191; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_193 = 6'h29 == value ? 32'h0 : _GEN_192; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_194 = 6'h2a == value ? 32'h0 : _GEN_193; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_195 = 6'h2b == value ? 32'h0 : _GEN_194; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_196 = 6'h2c == value ? 32'h0 : _GEN_195; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_197 = 6'h2d == value ? 32'h1 : _GEN_196; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_198 = 6'h2e == value ? 32'h0 : _GEN_197; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_199 = 6'h2f == value ? 32'h0 : _GEN_198; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_200 = 6'h30 == value ? 32'h1 : _GEN_199; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_201 = 6'h31 == value ? 32'h0 : _GEN_200; // @[ALUTests.scala 34:17:@1463.4]
  assign _T_1678 = _T_1665 ? _GEN_201 : _T_1677; // @[ALUTests.scala 34:17:@1463.4]
  assign _GEN_203 = 6'h1 == value ? 32'h0 : 32'h1; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_204 = 6'h2 == value ? 32'h1 : _GEN_203; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_205 = 6'h3 == value ? 32'h0 : _GEN_204; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_206 = 6'h4 == value ? 32'h1 : _GEN_205; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_207 = 6'h5 == value ? 32'h0 : _GEN_206; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_208 = 6'h6 == value ? 32'h0 : _GEN_207; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_209 = 6'h7 == value ? 32'h0 : _GEN_208; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_210 = 6'h8 == value ? 32'h1 : _GEN_209; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_211 = 6'h9 == value ? 32'h0 : _GEN_210; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_212 = 6'ha == value ? 32'h1 : _GEN_211; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_213 = 6'hb == value ? 32'h1 : _GEN_212; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_214 = 6'hc == value ? 32'h1 : _GEN_213; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_215 = 6'hd == value ? 32'h1 : _GEN_214; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_216 = 6'he == value ? 32'h0 : _GEN_215; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_217 = 6'hf == value ? 32'h0 : _GEN_216; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_218 = 6'h10 == value ? 32'h0 : _GEN_217; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_219 = 6'h11 == value ? 32'h1 : _GEN_218; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_220 = 6'h12 == value ? 32'h1 : _GEN_219; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_221 = 6'h13 == value ? 32'h1 : _GEN_220; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_222 = 6'h14 == value ? 32'h0 : _GEN_221; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_223 = 6'h15 == value ? 32'h0 : _GEN_222; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_224 = 6'h16 == value ? 32'h1 : _GEN_223; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_225 = 6'h17 == value ? 32'h1 : _GEN_224; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_226 = 6'h18 == value ? 32'h1 : _GEN_225; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_227 = 6'h19 == value ? 32'h0 : _GEN_226; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_228 = 6'h1a == value ? 32'h0 : _GEN_227; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_229 = 6'h1b == value ? 32'h1 : _GEN_228; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_230 = 6'h1c == value ? 32'h0 : _GEN_229; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_231 = 6'h1d == value ? 32'h0 : _GEN_230; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_232 = 6'h1e == value ? 32'h1 : _GEN_231; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_233 = 6'h1f == value ? 32'h1 : _GEN_232; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_234 = 6'h20 == value ? 32'h1 : _GEN_233; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_235 = 6'h21 == value ? 32'h1 : _GEN_234; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_236 = 6'h22 == value ? 32'h1 : _GEN_235; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_237 = 6'h23 == value ? 32'h0 : _GEN_236; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_238 = 6'h24 == value ? 32'h0 : _GEN_237; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_239 = 6'h25 == value ? 32'h0 : _GEN_238; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_240 = 6'h26 == value ? 32'h1 : _GEN_239; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_241 = 6'h27 == value ? 32'h0 : _GEN_240; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_242 = 6'h28 == value ? 32'h0 : _GEN_241; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_243 = 6'h29 == value ? 32'h1 : _GEN_242; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_244 = 6'h2a == value ? 32'h1 : _GEN_243; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_245 = 6'h2b == value ? 32'h0 : _GEN_244; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_246 = 6'h2c == value ? 32'h0 : _GEN_245; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_247 = 6'h2d == value ? 32'h0 : _GEN_246; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_248 = 6'h2e == value ? 32'h1 : _GEN_247; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_249 = 6'h2f == value ? 32'h0 : _GEN_248; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_250 = 6'h30 == value ? 32'h1 : _GEN_249; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_251 = 6'h31 == value ? 32'h0 : _GEN_250; // @[ALUTests.scala 33:17:@1464.4]
  assign _T_1679 = _T_1663 ? _GEN_251 : _T_1678; // @[ALUTests.scala 33:17:@1464.4]
  assign _GEN_253 = 6'h1 == value ? 32'hdcb6c7cd : 32'h50099a1c; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_254 = 6'h2 == value ? 32'h91dea927 : _GEN_253; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_255 = 6'h3 == value ? 32'h9cb48f7b : _GEN_254; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_256 = 6'h4 == value ? 32'h7b685ff7 : _GEN_255; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_257 = 6'h5 == value ? 32'hb0469759 : _GEN_256; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_258 = 6'h6 == value ? 32'hc2f739cd : _GEN_257; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_259 = 6'h7 == value ? 32'hddf254be : _GEN_258; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_260 = 6'h8 == value ? 32'h4ea4034 : _GEN_259; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_261 = 6'h9 == value ? 32'hbe03e3b8 : _GEN_260; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_262 = 6'ha == value ? 32'hb45aecba : _GEN_261; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_263 = 6'hb == value ? 32'ha3474102 : _GEN_262; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_264 = 6'hc == value ? 32'h300f5152 : _GEN_263; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_265 = 6'hd == value ? 32'h87e24ae : _GEN_264; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_266 = 6'he == value ? 32'h127d9d08 : _GEN_265; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_267 = 6'hf == value ? 32'hcf760c09 : _GEN_266; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_268 = 6'h10 == value ? 32'h9cfaf04 : _GEN_267; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_269 = 6'h11 == value ? 32'hbf557bd5 : _GEN_268; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_270 = 6'h12 == value ? 32'h1d3a5e78 : _GEN_269; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_271 = 6'h13 == value ? 32'hac31750 : _GEN_270; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_272 = 6'h14 == value ? 32'he0db3fcd : _GEN_271; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_273 = 6'h15 == value ? 32'h360feafc : _GEN_272; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_274 = 6'h16 == value ? 32'h20352b9e : _GEN_273; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_275 = 6'h17 == value ? 32'h4ea9b53e : _GEN_274; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_276 = 6'h18 == value ? 32'h5e1cb5d2 : _GEN_275; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_277 = 6'h19 == value ? 32'ha42c63b3 : _GEN_276; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_278 = 6'h1a == value ? 32'h75eb4d9f : _GEN_277; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_279 = 6'h1b == value ? 32'h29e729ff : _GEN_278; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_280 = 6'h1c == value ? 32'ha04bb81f : _GEN_279; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_281 = 6'h1d == value ? 32'h126dcd98 : _GEN_280; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_282 = 6'h1e == value ? 32'hc55bc572 : _GEN_281; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_283 = 6'h1f == value ? 32'hd63942d4 : _GEN_282; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_284 = 6'h20 == value ? 32'h2a505105 : _GEN_283; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_285 = 6'h21 == value ? 32'h74950fd7 : _GEN_284; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_286 = 6'h22 == value ? 32'hcb61cdc8 : _GEN_285; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_287 = 6'h23 == value ? 32'h82f8ab58 : _GEN_286; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_288 = 6'h24 == value ? 32'h82fc68c0 : _GEN_287; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_289 = 6'h25 == value ? 32'hfdf8a42b : _GEN_288; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_290 = 6'h26 == value ? 32'h6f6bb7dc : _GEN_289; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_291 = 6'h27 == value ? 32'hc476da0c : _GEN_290; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_292 = 6'h28 == value ? 32'h2ec9316f : _GEN_291; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_293 = 6'h29 == value ? 32'ha45ddc5e : _GEN_292; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_294 = 6'h2a == value ? 32'hcb3fbd57 : _GEN_293; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_295 = 6'h2b == value ? 32'h2cdb8fdb : _GEN_294; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_296 = 6'h2c == value ? 32'h3ba52ef : _GEN_295; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_297 = 6'h2d == value ? 32'haa6dc03d : _GEN_296; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_298 = 6'h2e == value ? 32'h834f41bb : _GEN_297; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_299 = 6'h2f == value ? 32'h69c01cb5 : _GEN_298; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_300 = 6'h30 == value ? 32'h12e81440 : _GEN_299; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_301 = 6'h31 == value ? 32'h2c951562 : _GEN_300; // @[ALUTests.scala 32:17:@1465.4]
  assign _T_1680 = _T_1661 ? _GEN_301 : _T_1679; // @[ALUTests.scala 32:17:@1465.4]
  assign _GEN_303 = 6'h1 == value ? 32'hffb7d7cd : 32'hd489bfbd; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_304 = 6'h2 == value ? 32'hbbdefdbf : _GEN_303; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_305 = 6'h3 == value ? 32'h9db5cf7b : _GEN_304; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_306 = 6'h4 == value ? 32'h7f6bfff7 : _GEN_305; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_307 = 6'h5 == value ? 32'hb4e7975b : _GEN_306; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_308 = 6'h6 == value ? 32'hcaf7fbff : _GEN_307; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_309 = 6'h7 == value ? 32'hddfbd6ff : _GEN_308; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_310 = 6'h8 == value ? 32'heceae235 : _GEN_309; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_311 = 6'h9 == value ? 32'hfe67f7fe : _GEN_310; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_312 = 6'ha == value ? 32'hbf5fedbb : _GEN_311; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_313 = 6'hb == value ? 32'hab7fd3b3 : _GEN_312; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_314 = 6'hc == value ? 32'h70cf7756 : _GEN_313; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_315 = 6'hd == value ? 32'h7efe34ae : _GEN_314; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_316 = 6'he == value ? 32'h5f7dbfab : _GEN_315; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_317 = 6'hf == value ? 32'hdff69f9b : _GEN_316; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_318 = 6'h10 == value ? 32'hfdfafb5 : _GEN_317; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_319 = 6'h11 == value ? 32'hfff5fbfd : _GEN_318; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_320 = 6'h12 == value ? 32'h5d3f7efa : _GEN_319; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_321 = 6'h13 == value ? 32'heefb57fa : _GEN_320; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_322 = 6'h14 == value ? 32'he2ffbfff : _GEN_321; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_323 = 6'h15 == value ? 32'hb6affefc : _GEN_322; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_324 = 6'h16 == value ? 32'h327dabff : _GEN_323; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_325 = 6'h17 == value ? 32'hefadfdbe : _GEN_324; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_326 = 6'h18 == value ? 32'hfe7cbfde : _GEN_325; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_327 = 6'h19 == value ? 32'hf76e73f3 : _GEN_326; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_328 = 6'h1a == value ? 32'h7def7fff : _GEN_327; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_329 = 6'h1b == value ? 32'hf9ff6bff : _GEN_328; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_330 = 6'h1c == value ? 32'hbd5bfd1f : _GEN_329; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_331 = 6'h1d == value ? 32'h93fdcfbc : _GEN_330; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_332 = 6'h1e == value ? 32'hddffedf3 : _GEN_331; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_333 = 6'h1f == value ? 32'hde7fe6ff : _GEN_332; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_334 = 6'h20 == value ? 32'hba59d5a7 : _GEN_333; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_335 = 6'h21 == value ? 32'hfed5aff7 : _GEN_334; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_336 = 6'h22 == value ? 32'hef79cdde : _GEN_335; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_337 = 6'h23 == value ? 32'haffbeb5c : _GEN_336; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_338 = 6'h24 == value ? 32'hf3fc7fc7 : _GEN_337; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_339 = 6'h25 == value ? 32'hfdfced3f : _GEN_338; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_340 = 6'h26 == value ? 32'heffbf7dd : _GEN_339; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_341 = 6'h27 == value ? 32'hc7f7fe2e : _GEN_340; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_342 = 6'h28 == value ? 32'hafcff77f : _GEN_341; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_343 = 6'h29 == value ? 32'hac7ddddf : _GEN_342; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_344 = 6'h2a == value ? 32'hebbffff7 : _GEN_343; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_345 = 6'h2b == value ? 32'hadff8fdb : _GEN_344; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_346 = 6'h2c == value ? 32'h23ba7bef : _GEN_345; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_347 = 6'h2d == value ? 32'hbe6deffd : _GEN_346; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_348 = 6'h2e == value ? 32'ha7dff3fb : _GEN_347; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_349 = 6'h2f == value ? 32'hefc95eb7 : _GEN_348; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_350 = 6'h30 == value ? 32'hbaecffcb : _GEN_349; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_351 = 6'h31 == value ? 32'h6ef5d7f6 : _GEN_350; // @[ALUTests.scala 31:17:@1466.4]
  assign _T_1681 = _T_1659 ? _GEN_351 : _T_1680; // @[ALUTests.scala 31:17:@1466.4]
  assign _GEN_353 = 6'h1 == value ? 32'h23011000 : 32'h848025a1; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_354 = 6'h2 == value ? 32'h2a005498 : _GEN_353; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_355 = 6'h3 == value ? 32'h1014000 : _GEN_354; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_356 = 6'h4 == value ? 32'h403a000 : _GEN_355; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_357 = 6'h5 == value ? 32'h4a10002 : _GEN_356; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_358 = 6'h6 == value ? 32'h800c232 : _GEN_357; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_359 = 6'h7 == value ? 32'h98241 : _GEN_358; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_360 = 6'h8 == value ? 32'he800a201 : _GEN_359; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_361 = 6'h9 == value ? 32'h40641446 : _GEN_360; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_362 = 6'ha == value ? 32'hb050101 : _GEN_361; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_363 = 6'hb == value ? 32'h83892b1 : _GEN_362; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_364 = 6'hc == value ? 32'h40c02604 : _GEN_363; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_365 = 6'hd == value ? 32'h76801000 : _GEN_364; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_366 = 6'he == value ? 32'h4d0022a3 : _GEN_365; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_367 = 6'hf == value ? 32'h10809392 : _GEN_366; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_368 = 6'h10 == value ? 32'h61000b1 : _GEN_367; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_369 = 6'h11 == value ? 32'h40a08028 : _GEN_368; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_370 = 6'h12 == value ? 32'h40052082 : _GEN_369; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_371 = 6'h13 == value ? 32'he43840aa : _GEN_370; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_372 = 6'h14 == value ? 32'h2248032 : _GEN_371; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_373 = 6'h15 == value ? 32'h80a01400 : _GEN_372; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_374 = 6'h16 == value ? 32'h12488061 : _GEN_373; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_375 = 6'h17 == value ? 32'ha1044880 : _GEN_374; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_376 = 6'h18 == value ? 32'ha0600a0c : _GEN_375; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_377 = 6'h19 == value ? 32'h53421040 : _GEN_376; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_378 = 6'h1a == value ? 32'h8043260 : _GEN_377; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_379 = 6'h1b == value ? 32'hd0184200 : _GEN_378; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_380 = 6'h1c == value ? 32'h1d104500 : _GEN_379; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_381 = 6'h1d == value ? 32'h81900224 : _GEN_380; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_382 = 6'h1e == value ? 32'h18a42881 : _GEN_381; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_383 = 6'h1f == value ? 32'h846a42b : _GEN_382; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_384 = 6'h20 == value ? 32'h900984a2 : _GEN_383; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_385 = 6'h21 == value ? 32'h8a40a020 : _GEN_384; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_386 = 6'h22 == value ? 32'h24180016 : _GEN_385; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_387 = 6'h23 == value ? 32'h2d034004 : _GEN_386; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_388 = 6'h24 == value ? 32'h71001707 : _GEN_387; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_389 = 6'h25 == value ? 32'h44914 : _GEN_388; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_390 = 6'h26 == value ? 32'h80904001 : _GEN_389; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_391 = 6'h27 == value ? 32'h3812422 : _GEN_390; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_392 = 6'h28 == value ? 32'h8106c610 : _GEN_391; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_393 = 6'h29 == value ? 32'h8200181 : _GEN_392; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_394 = 6'h2a == value ? 32'h208042a0 : _GEN_393; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_395 = 6'h2b == value ? 32'h81240000 : _GEN_394; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_396 = 6'h2c == value ? 32'h20002900 : _GEN_395; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_397 = 6'h2d == value ? 32'h14002fc0 : _GEN_396; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_398 = 6'h2e == value ? 32'h2490b240 : _GEN_397; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_399 = 6'h2f == value ? 32'h86094202 : _GEN_398; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_400 = 6'h30 == value ? 32'ha804eb8b : _GEN_399; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_401 = 6'h31 == value ? 32'h4260c294 : _GEN_400; // @[ALUTests.scala 30:17:@1467.4]
  assign _T_1682 = _T_1657 ? _GEN_401 : _T_1681; // @[ALUTests.scala 30:17:@1467.4]
  assign _GEN_403 = 6'h1 == value ? 32'hdb693b43 : 32'hcff779ec; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_404 = 6'h2 == value ? 32'h6ede68e5 : _GEN_403; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_405 = 6'h3 == value ? 32'h9c938165 : _GEN_404; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_406 = 6'h4 == value ? 32'hf567d7ef : _GEN_405; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_407 = 6'h5 == value ? 32'hb03e6ab7 : _GEN_406; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_408 = 6'h6 == value ? 32'hbdccc7c3 : _GEN_407; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_409 = 6'h7 == value ? 32'hd232339a : _GEN_408; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_410 = 6'h8 == value ? 32'hfbd6400c : _GEN_409; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_411 = 6'h9 == value ? 32'h4e01dca8 : _GEN_410; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_412 = 6'ha == value ? 32'h6bd9946a : _GEN_411; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_413 = 6'hb == value ? 32'h5f393f02 : _GEN_412; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_414 = 6'hc == value ? 32'hf002d0ae : _GEN_413; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_415 = 6'hd == value ? 32'hf7ae236a : _GEN_414; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_416 = 6'he == value ? 32'he356b08 : _GEN_415; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_417 = 6'hf == value ? 32'hb949f3f9 : _GEN_416; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_418 = 6'h10 == value ? 32'h74b58fc : _GEN_417; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_419 = 6'h11 == value ? 32'h9b54c635 : _GEN_418; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_420 = 6'h12 == value ? 32'heae5d1b8 : _GEN_419; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_421 = 6'h13 == value ? 32'hf6411130 : _GEN_420; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_422 = 6'h14 == value ? 32'h60c4e6bb : _GEN_421; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_423 = 6'h15 == value ? 32'h9f6e98c : _GEN_422; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_424 = 6'h16 == value ? 32'hdfcb2962 : _GEN_423; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_425 = 6'h17 == value ? 32'hcea7930e : _GEN_424; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_426 = 6'h18 == value ? 32'hd6145232 : _GEN_425; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_427 = 6'h19 == value ? 32'ha3e41d93 : _GEN_426; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_428 = 6'h1a == value ? 32'h74e8cc9d : _GEN_427; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_429 = 6'h1b == value ? 32'he8a51911 : _GEN_428; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_430 = 6'h1c == value ? 32'h6037a7ff : _GEN_429; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_431 = 6'h1d == value ? 32'h121bb278 : _GEN_430; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_432 = 6'h1e == value ? 32'h45243c8e : _GEN_431; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_433 = 6'h1f == value ? 32'hd237412c : _GEN_432; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_434 = 6'h20 == value ? 32'hd9b05105 : _GEN_433; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_435 = 6'h21 == value ? 32'hd492f2cd : _GEN_434; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_436 = 6'h22 == value ? 32'hbb1e3bc8 : _GEN_435; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_437 = 6'h23 == value ? 32'h7e475928 : _GEN_436; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_438 = 6'h24 == value ? 32'h829bd840 : _GEN_437; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_439 = 6'h25 == value ? 32'h6d08a3eb : _GEN_438; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_440 = 6'h26 == value ? 32'heb16b72c : _GEN_439; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_441 = 6'h27 == value ? 32'hbc6dc604 : _GEN_440; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_442 = 6'h28 == value ? 32'h1a472ead : _GEN_441; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_443 = 6'h29 == value ? 32'h64342c4e : _GEN_442; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_444 = 6'h2a == value ? 32'hc4fa5cc9 : _GEN_443; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_445 = 6'h2b == value ? 32'h14c88157 : _GEN_444; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_446 = 6'h2c == value ? 32'h2a64d25 : _GEN_445; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_447 = 6'h2d == value ? 32'h59a4bffd : _GEN_446; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_448 = 6'h2e == value ? 32'h80c6c0bb : _GEN_447; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_449 = 6'h2f == value ? 32'h26400cab : _GEN_448; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_450 = 6'h30 == value ? 32'hf2d81440 : _GEN_449; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_451 = 6'h31 == value ? 32'h238af2e2 : _GEN_450; // @[ALUTests.scala 29:17:@1468.4]
  assign _T_1683 = _T_1655 ? _GEN_451 : _T_1682; // @[ALUTests.scala 29:17:@1468.4]
  assign _GEN_453 = 6'h1 == value ? 32'h22b8e7cd : 32'h5909e55e; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_454 = 6'h2 == value ? 32'he5df5257 : _GEN_453; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_455 = 6'h3 == value ? 32'h9eb70f7b : _GEN_454; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_456 = 6'h4 == value ? 32'h836f9ff7 : _GEN_455; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_457 = 6'h5 == value ? 32'hb988975d : _GEN_456; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_458 = 6'h6 == value ? 32'hd2f8be31 : _GEN_457; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_459 = 6'h7 == value ? 32'hde055940 : _GEN_458; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_460 = 6'h8 == value ? 32'hd4eb8436 : _GEN_459; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_461 = 6'h9 == value ? 32'h3ecc0c44 : _GEN_460; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_462 = 6'ha == value ? 32'hca64eebc : _GEN_461; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_463 = 6'hb == value ? 32'hb3b86664 : _GEN_462; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_464 = 6'hc == value ? 32'hb18f9d5a : _GEN_463; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_465 = 6'hd == value ? 32'hf57e44ae : _GEN_464; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_466 = 6'he == value ? 32'hac7de24e : _GEN_465; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_467 = 6'hf == value ? 32'hf077332d : _GEN_466; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_468 = 6'h10 == value ? 32'h15efb066 : _GEN_467; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_469 = 6'h11 == value ? 32'h40967c25 : _GEN_468; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_470 = 6'h12 == value ? 32'h9d449f7c : _GEN_469; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_471 = 6'h13 == value ? 32'hd33398a4 : _GEN_470; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_472 = 6'h14 == value ? 32'he5244031 : _GEN_471; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_473 = 6'h15 == value ? 32'h375012fc : _GEN_472; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_474 = 6'h16 == value ? 32'h44c62c60 : _GEN_473; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_475 = 6'h17 == value ? 32'h90b2463e : _GEN_474; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_476 = 6'h18 == value ? 32'h9edcc9ea : _GEN_475; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_477 = 6'h19 == value ? 32'h4ab08433 : _GEN_476; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_478 = 6'h1a == value ? 32'h85f3b25f : _GEN_477; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_479 = 6'h1b == value ? 32'hca17adff : _GEN_478; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_480 = 6'h1c == value ? 32'hda6c421f : _GEN_479; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_481 = 6'h1d == value ? 32'h158dd1e0 : _GEN_480; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_482 = 6'h1e == value ? 32'hf6a41674 : _GEN_481; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_483 = 6'h1f == value ? 32'he6c68b2a : _GEN_482; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_484 = 6'h20 == value ? 32'h4a635a49 : _GEN_483; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_485 = 6'h21 == value ? 32'h89165017 : _GEN_484; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_486 = 6'h22 == value ? 32'h1391cdf4 : _GEN_485; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_487 = 6'h23 == value ? 32'hdcff2b60 : _GEN_486; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_488 = 6'h24 == value ? 32'h64fc96ce : _GEN_487; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_489 = 6'h25 == value ? 32'hfe013653 : _GEN_488; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_490 = 6'h26 == value ? 32'h708c37de : _GEN_489; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_491 = 6'h27 == value ? 32'hcb792250 : _GEN_490; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_492 = 6'h28 == value ? 32'h30d6bd8f : _GEN_491; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_493 = 6'h29 == value ? 32'hb49ddf60 : _GEN_492; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_494 = 6'h2a == value ? 32'hc404297 : _GEN_493; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_495 = 6'h2b == value ? 32'h2f238fdb : _GEN_494; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_496 = 6'h2c == value ? 32'h43baa4ef : _GEN_495; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_497 = 6'h2d == value ? 32'hd26e1fbd : _GEN_496; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_498 = 6'h2e == value ? 32'hcc70a63b : _GEN_497; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_499 = 6'h2f == value ? 32'h75d2a0b9 : _GEN_498; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_500 = 6'h30 == value ? 32'h62f1eb56 : _GEN_499; // @[ALUTests.scala 28:17:@1469.4]
  assign _GEN_501 = 6'h31 == value ? 32'hb1569a8a : _GEN_500; // @[ALUTests.scala 28:17:@1469.4]
  assign _T_1684 = _T_1653 ? _GEN_501 : _T_1683; // @[ALUTests.scala 28:17:@1469.4]
  assign _T_1685 = dut_io_alu_op[0]; // @[ALUTests.scala 39:31:@1470.4]
  assign _T_1688 = _T_1685 ? _GEN_451 : _GEN_501; // @[ALUTests.scala 39:17:@1471.4]
  assign _GEN_503 = 6'h1 == value ? 32'h693ef17 : 32'hefe57db7; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_504 = 6'h2 == value ? 32'hb7727a6f : _GEN_503; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_505 = 6'h3 == value ? 32'haf120267 : _GEN_504; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_506 = 6'h4 == value ? 32'h4ecc00e3 : _GEN_505; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_507 = 6'h5 == value ? 32'he84191e3 : _GEN_506; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_508 = 6'h6 == value ? 32'h194acfe3 : _GEN_507; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_509 = 6'h7 == value ? 32'hb834d363 : _GEN_508; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_510 = 6'h8 == value ? 32'h3bfeebe3 : _GEN_509; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_511 = 6'h9 == value ? 32'h630af363 : _GEN_510; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_512 = 6'ha == value ? 32'h18ec0483 : _GEN_511; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_513 = 6'hb == value ? 32'hcfc9603 : _GEN_512; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_514 = 6'hc == value ? 32'hbe742b83 : _GEN_513; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_515 = 6'hd == value ? 32'h3352c283 : _GEN_514; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_516 = 6'he == value ? 32'h5cc25c83 : _GEN_515; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_517 = 6'hf == value ? 32'h8af40923 : _GEN_516; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_518 = 6'h10 == value ? 32'hb6d81fa3 : _GEN_517; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_519 = 6'h11 == value ? 32'hc903aba3 : _GEN_518; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_520 = 6'h12 == value ? 32'hfd2e8913 : _GEN_519; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_521 = 6'h13 == value ? 32'hbfdad93 : _GEN_520; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_522 = 6'h14 == value ? 32'h37fbb093 : _GEN_521; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_523 = 6'h15 == value ? 32'hee814093 : _GEN_522; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_524 = 6'h16 == value ? 32'hd05eea13 : _GEN_523; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_525 = 6'h17 == value ? 32'h388cf313 : _GEN_524; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_526 = 6'h18 == value ? 32'hfd1293 : _GEN_525; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_527 = 6'h19 == value ? 32'h162df93 : _GEN_526; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_528 = 6'h1a == value ? 32'h41435713 : _GEN_527; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_529 = 6'h1b == value ? 32'h4a8eb3 : _GEN_528; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_530 = 6'h1c == value ? 32'h41d90c33 : _GEN_529; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_531 = 6'h1d == value ? 32'h7e97b3 : _GEN_530; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_532 = 6'h1e == value ? 32'h32af33 : _GEN_531; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_533 = 6'h1f == value ? 32'h863833 : _GEN_532; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_534 = 6'h20 == value ? 32'hc4c133 : _GEN_533; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_535 = 6'h21 == value ? 32'h121d633 : _GEN_534; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_536 = 6'h22 == value ? 32'h40ecdf33 : _GEN_535; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_537 = 6'h23 == value ? 32'h326d33 : _GEN_536; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_538 = 6'h24 == value ? 32'h16df6b3 : _GEN_537; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_539 = 6'h25 == value ? 32'hff0000f : _GEN_538; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_540 = 6'h26 == value ? 32'h100f : _GEN_539; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_541 = 6'h27 == value ? 32'hc82c13f3 : _GEN_540; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_542 = 6'h28 == value ? 32'h34142673 : _GEN_541; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_543 = 6'h29 == value ? 32'h344c35f3 : _GEN_542; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_544 = 6'h2a == value ? 32'h780656f3 : _GEN_543; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_545 = 6'h2b == value ? 32'h701a6173 : _GEN_544; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_546 = 6'h2c == value ? 32'hf01d76f3 : _GEN_545; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_547 = 6'h2d == value ? 32'h73 : _GEN_546; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_548 = 6'h2e == value ? 32'h100073 : _GEN_547; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_549 = 6'h2f == value ? 32'h10000073 : _GEN_548; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_550 = 6'h30 == value ? 32'h13 : _GEN_549; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_551 = 6'h31 == value ? 32'h1e2b73b3 : _GEN_550; // @[ALUTests.scala 41:16:@1523.4]
  assign _GEN_553 = 6'h1 == value ? 32'h7f111188 : 32'h9480afa5; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_554 = 6'h2 == value ? 32'haa5edd9e : _GEN_553; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_555 = 6'h3 == value ? 32'h1da54870 : _GEN_554; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_556 = 6'h4 == value ? 32'h3c6bbbf3 : _GEN_555; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_557 = 6'h5 == value ? 32'h34e3810a : _GEN_556; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_558 = 6'h6 == value ? 32'h4862c2fa : _GEN_557; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_559 = 6'h7 == value ? 32'h581bc66d : _GEN_558; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_560 = 6'h8 == value ? 32'he860e221 : _GEN_559; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_561 = 6'h9 == value ? 32'h4666f476 : _GEN_560; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_562 = 6'ha == value ? 32'h9b1f4193 : _GEN_561; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_563 = 6'hb == value ? 32'h8978d2b3 : _GEN_562; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_564 = 6'hc == value ? 32'h50c93704 : _GEN_563; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_565 = 6'hd == value ? 32'h7696340c : _GEN_564; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_566 = 6'he == value ? 32'h5d59a6ab : _GEN_565; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_567 = 6'hf == value ? 32'h54e09393 : _GEN_566; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_568 = 6'h10 == value ? 32'he9d84b1 : _GEN_567; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_569 = 6'h11 == value ? 32'hedf5a12d : _GEN_568; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_570 = 6'h12 == value ? 32'h4415389a : _GEN_569; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_571 = 6'h13 == value ? 32'he4ba54ea : _GEN_570; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_572 = 6'h14 == value ? 32'h22f49376 : _GEN_571; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_573 = 6'h15 == value ? 32'ha0a37e44 : _GEN_572; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_574 = 6'h16 == value ? 32'h1248aae1 : _GEN_573; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_575 = 6'h17 == value ? 32'hafaceca6 : _GEN_574; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_576 = 6'h18 == value ? 32'hba788e0e : _GEN_575; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_577 = 6'h19 == value ? 32'h774a50e3 : _GEN_576; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_578 = 6'h1a == value ? 32'h7d6e3f7e : _GEN_577; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_579 = 6'h1b == value ? 32'hd95e6388 : _GEN_578; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_580 = 6'h1c == value ? 32'h1d51f50f : _GEN_579; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_581 = 6'h1d == value ? 32'h93d4c22c : _GEN_580; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_582 = 6'h1e == value ? 32'h9de42981 : _GEN_581; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_583 = 6'h1f == value ? 32'hdc7ee62b : _GEN_582; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_584 = 6'h20 == value ? 32'h9209d5a7 : _GEN_583; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_585 = 6'h21 == value ? 32'haed4a172 : _GEN_584; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_586 = 6'h22 == value ? 32'he75804de : _GEN_585; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_587 = 6'h23 == value ? 32'h2da34244 : _GEN_586; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_588 = 6'h24 == value ? 32'h73cc3787 : _GEN_587; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_589 = 6'h25 == value ? 32'h3584ed1f : _GEN_588; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_590 = 6'h26 == value ? 32'hadd17785 : _GEN_589; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_591 = 6'h27 == value ? 32'h43f3742a : _GEN_590; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_592 = 6'h28 == value ? 32'ha58ef61e : _GEN_591; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_593 = 6'h29 == value ? 32'h8c6905d7 : _GEN_592; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_594 = 6'h2a == value ? 32'he89d4fb0 : _GEN_593; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_595 = 6'h2b == value ? 32'ha1f60899 : _GEN_594; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_596 = 6'h2c == value ? 32'h2330790a : _GEN_595; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_597 = 6'h2d == value ? 32'h16096fdd : _GEN_596; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_598 = 6'h2e == value ? 32'ha69bb37b : _GEN_597; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_599 = 6'h2f == value ? 32'hce0956b2 : _GEN_598; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_600 = 6'h30 == value ? 32'haae4ffcb : _GEN_599; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_601 = 6'h31 == value ? 32'h6a70c6b6 : _GEN_600; // @[ALUTests.scala 43:12:@1576.4]
  assign _GEN_603 = 6'h1 == value ? 32'ha3a7d645 : 32'hc48935b9; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_604 = 6'h2 == value ? 32'h3b8074b9 : _GEN_603; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_605 = 6'h3 == value ? 32'h8111c70b : _GEN_604; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_606 = 6'h4 == value ? 32'h4703e404 : _GEN_605; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_607 = 6'h5 == value ? 32'h84a51653 : _GEN_606; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_608 = 6'h6 == value ? 32'h8a95fb37 : _GEN_607; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_609 = 6'h7 == value ? 32'h85e992d3 : _GEN_608; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_610 = 6'h8 == value ? 32'hec8aa215 : _GEN_609; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_611 = 6'h9 == value ? 32'hf86517ce : _GEN_610; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_612 = 6'ha == value ? 32'h2f45ad29 : _GEN_611; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_613 = 6'hb == value ? 32'h2a3f93b1 : _GEN_612; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_614 = 6'hc == value ? 32'h60c66656 : _GEN_613; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_615 = 6'hd == value ? 32'h7ee810a2 : _GEN_614; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_616 = 6'he == value ? 32'h4f243ba3 : _GEN_615; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_617 = 6'hf == value ? 32'h9b969f9a : _GEN_616; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_618 = 6'h10 == value ? 32'h7522bb5 : _GEN_617; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_619 = 6'h11 == value ? 32'h52a0daf8 : _GEN_618; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_620 = 6'h12 == value ? 32'h592f66e2 : _GEN_619; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_621 = 6'h13 == value ? 32'hee7943ba : _GEN_620; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_622 = 6'h14 == value ? 32'hc22facbb : _GEN_621; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_623 = 6'h15 == value ? 32'h96ac94b8 : _GEN_622; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_624 = 6'h16 == value ? 32'h327d817f : _GEN_623; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_625 = 6'h17 == value ? 32'he1055998 : _GEN_624; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_626 = 6'h18 == value ? 32'he4643bdc : _GEN_625; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_627 = 6'h19 == value ? 32'hd3663350 : _GEN_626; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_628 = 6'h1a == value ? 32'h88572e1 : _GEN_627; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_629 = 6'h1b == value ? 32'hf0b94a77 : _GEN_628; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_630 = 6'h1c == value ? 32'hbd1a4d10 : _GEN_629; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_631 = 6'h1d == value ? 32'h81b90fb4 : _GEN_630; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_632 = 6'h1e == value ? 32'h58bfecf3 : _GEN_631; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_633 = 6'h1f == value ? 32'ha47a4ff : _GEN_632; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_634 = 6'h20 == value ? 32'hb85984a2 : _GEN_633; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_635 = 6'h21 == value ? 32'hda41aea5 : _GEN_634; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_636 = 6'h22 == value ? 32'h2c39c916 : _GEN_635; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_637 = 6'h23 == value ? 32'haf5be91c : _GEN_636; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_638 = 6'h24 == value ? 32'hf1305f47 : _GEN_637; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_639 = 6'h25 == value ? 32'hc87c4934 : _GEN_638; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_640 = 6'h26 == value ? 32'hc2bac059 : _GEN_639; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_641 = 6'h27 == value ? 32'h8785ae26 : _GEN_640; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_642 = 6'h28 == value ? 32'h8b47c771 : _GEN_641; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_643 = 6'h29 == value ? 32'h2834d989 : _GEN_642; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_644 = 6'h2a == value ? 32'h23a2f2e7 : _GEN_643; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_645 = 6'h2b == value ? 32'h8d2d8742 : _GEN_644; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_646 = 6'h2c == value ? 32'h208a2be5 : _GEN_645; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_647 = 6'h2d == value ? 32'hbc64afe0 : _GEN_646; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_648 = 6'h2e == value ? 32'h25d4f2c0 : _GEN_647; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_649 = 6'h2f == value ? 32'ha7c94a07 : _GEN_648; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_650 = 6'h30 == value ? 32'hb80ceb8b : _GEN_649; // @[ALUTests.scala 44:12:@1628.4]
  assign _GEN_651 = 6'h31 == value ? 32'h46e5d3d4 : _GEN_650; // @[ALUTests.scala 44:12:@1628.4]
  assign _T_1959 = reset == 1'h0; // @[ALUTests.scala 46:20:@1631.6]
  assign _T_1963 = dut_io_out == _T_1684; // @[ALUTests.scala 47:21:@1641.4]
  assign _T_1965 = _T_1963 | reset; // @[ALUTests.scala 47:9:@1643.4]
  assign _T_1967 = _T_1965 == 1'h0; // @[ALUTests.scala 47:9:@1644.4]
  assign _T_1968 = dut_io_sum == _T_1688; // @[ALUTests.scala 48:21:@1649.4]
  assign _T_1970 = _T_1968 | reset; // @[ALUTests.scala 48:9:@1651.4]
  assign _T_1972 = _T_1970 == 1'h0; // @[ALUTests.scala 48:9:@1652.4]
  assign dut_io_A = _GEN_601;
  assign dut_io_B = _GEN_651;
  assign dut_io_alu_op = ctrl_io_alu_op;
  assign ctrl_io_inst = _GEN_551;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  value = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      value <= 6'h0;
    end else begin
      if (done) begin
        value <= 6'h0;
      end else begin
        value <= _T_611;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (done & _T_1959) begin
          $finish; // @[ALUTests.scala 46:20:@1633.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (done & _T_1959) begin
          $finish; // @[ALUTests.scala 46:28:@1638.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1967) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ALUTests.scala:47 assert(dut.io.out === out._1)\n"); // @[ALUTests.scala 47:9:@1646.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1967) begin
          $fatal; // @[ALUTests.scala 47:9:@1647.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1972) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ALUTests.scala:48 assert(dut.io.sum === out._2)\n"); // @[ALUTests.scala 48:9:@1654.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1972) begin
          $fatal; // @[ALUTests.scala 48:9:@1655.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1959) begin
          $fwrite(32'h80000002,"Counter: %d, OP: 0x%h, A: 0x%h, B: 0x%h, OUT: 0x%h ?= 0x%h, SUM: 0x%h ?= 0x%h\n",value,dut_io_alu_op,dut_io_A,dut_io_B,dut_io_out,_T_1684,dut_io_sum,_T_1688); // @[ALUTests.scala 49:9:@1660.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
